module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [0:0] __in0,
  input logic [511:0] __in1,
  output logic [0:0] __out0,
  output logic [511:0] __out1);
  logic [6157:0] zll_pure_dispatch_in;
  logic [6155:0] zll_pure_dispatch4_in;
  logic [6155:0] zll_pure_dispatch5_in;
  logic [6155:0] zll_main_refold1_in;
  logic [5642:0] main_conn10_in;
  logic [5129:0] main_conn10_out;
  logic [5129:0] zll_main_ten11_in;
  logic [5129:0] zll_main_ten11_out;
  logic [5642:0] main_refold2_in;
  logic [6157:0] main_refold2_out;
  logic [6157:0] zll_pure_dispatch3_in;
  logic [512:0] main_refold_in;
  logic [5642:0] main_conn10_inR1;
  logic [5129:0] main_conn10_outR1;
  logic [5129:0] zll_main_ten11_inR1;
  logic [5129:0] zll_main_ten11_outR1;
  logic [5129:0] zll_main_out101_in;
  logic [512:0] zll_main_out101_out;
  logic [6157:0] zll_pure_dispatch1_in;
  logic [1025:0] zll_pure_dispatch2_in;
  logic [1025:0] zll_main_refold_in;
  logic [5642:0] main_conn10_inR2;
  logic [5129:0] main_conn10_outR2;
  logic [5129:0] zll_main_ten11_inR2;
  logic [5129:0] zll_main_ten11_outR2;
  logic [5642:0] main_refold2_inR1;
  logic [6157:0] main_refold2_outR1;
  logic [0:0] __continue;
  logic [5644:0] __resumption_tag;
  logic [5644:0] __resumption_tag_next;
  assign zll_pure_dispatch_in = {{__in0, __in1}, __resumption_tag};
  assign zll_pure_dispatch4_in = {zll_pure_dispatch_in[6157:5645], zll_pure_dispatch_in[5642:5130], zll_pure_dispatch_in[5129:0]};
  assign zll_pure_dispatch5_in = {zll_pure_dispatch4_in[5642:5130], zll_pure_dispatch4_in[6155:5643], zll_pure_dispatch4_in[5129:0]};
  assign zll_main_refold1_in = {zll_pure_dispatch5_in[6155:5643], zll_pure_dispatch5_in[5129:0], zll_pure_dispatch5_in[5642:5130]};
  assign main_conn10_in = {zll_main_refold1_in[5642:513], zll_main_refold1_in[6155:5643]};
  Main_conn10  inst (main_conn10_in[5642:513], main_conn10_in[512:0], main_conn10_out);
  assign zll_main_ten11_in = main_conn10_out;
  ZLL_Main_ten11  instR1 (zll_main_ten11_in[5129:0], zll_main_ten11_out);
  assign main_refold2_in = {zll_main_ten11_out, zll_main_refold1_in[512:0]};
  Main_refold2  instR2 (main_refold2_in[5642:513], main_refold2_in[512:0], main_refold2_out);
  assign zll_pure_dispatch3_in = {{__in0, __in1}, __resumption_tag};
  assign main_refold_in = zll_pure_dispatch3_in[6157:5645];
  assign main_conn10_inR1 = {{13'h140a{1'h0}}, main_refold_in[512:0]};
  Main_conn10  instR3 (main_conn10_inR1[5642:513], main_conn10_inR1[512:0], main_conn10_outR1);
  assign zll_main_ten11_inR1 = main_conn10_outR1;
  ZLL_Main_ten11  instR4 (zll_main_ten11_inR1[5129:0], zll_main_ten11_outR1);
  assign zll_main_out101_in = zll_main_ten11_outR1;
  ZLL_Main_out101  instR5 (zll_main_out101_in[5129:0], zll_main_out101_out);
  assign zll_pure_dispatch1_in = {{__in0, __in1}, __resumption_tag};
  assign zll_pure_dispatch2_in = {zll_pure_dispatch1_in[6157:5645], zll_pure_dispatch1_in[512:0]};
  assign zll_main_refold_in = {zll_pure_dispatch2_in[512:0], zll_pure_dispatch2_in[1025:513]};
  assign main_conn10_inR2 = {{13'h140a{1'h0}}, zll_main_refold_in[1025:513]};
  Main_conn10  instR6 (main_conn10_inR2[5642:513], main_conn10_inR2[512:0], main_conn10_outR2);
  assign zll_main_ten11_inR2 = main_conn10_outR2;
  ZLL_Main_ten11  instR7 (zll_main_ten11_inR2[5129:0], zll_main_ten11_outR2);
  assign main_refold2_inR1 = {zll_main_ten11_outR2, zll_main_refold_in[512:0]};
  Main_refold2  instR8 (main_refold2_inR1[5642:513], main_refold2_inR1[512:0], main_refold2_outR1);
  assign {__continue, __out0, __out1, __resumption_tag_next} = (zll_pure_dispatch1_in[5644:5643] == 2'h1) ? main_refold2_outR1 : ((zll_pure_dispatch3_in[5644:5643] == 2'h2) ? {zll_main_out101_out, {2'h1, {13'h140a{1'h0}}}, main_refold_in[512:0]} : main_refold2_out);
  initial __resumption_tag <= {1'h1, {13'h160c{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {1'h1, {13'h160c{1'h0}}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module ZLL_QuarterRound_quarterround39 (input logic [127:0] arg0,
  output logic [127:0] res);
  logic [127:0] zll_quarterround_quarterround34_in;
  logic [127:0] zll_quarterround_quarterround2_in;
  logic [63:0] binop_in;
  logic [31:0] zll_quarterround_quarterround28_in;
  logic [63:0] zll_quarterround_quarterround25_in;
  logic [31:0] zll_quarterround_quarterround25_out;
  logic [63:0] binop_inR1;
  logic [127:0] zll_quarterround_quarterround16_in;
  logic [63:0] binop_inR2;
  logic [31:0] zll_quarterround_quarterround4_in;
  logic [63:0] zll_quarterround_quarterround25_inR1;
  logic [31:0] zll_quarterround_quarterround25_outR1;
  logic [63:0] binop_inR3;
  logic [127:0] zll_quarterround_quarterround40_in;
  logic [63:0] binop_inR4;
  logic [31:0] zll_quarterround_quarterround12_in;
  logic [63:0] zll_quarterround_quarterround25_inR2;
  logic [31:0] zll_quarterround_quarterround25_outR2;
  logic [63:0] binop_inR5;
  logic [127:0] zll_quarterround_quarterround6_in;
  logic [63:0] binop_inR6;
  logic [31:0] zll_quarterround_quarterround17_in;
  logic [63:0] zll_quarterround_quarterround25_inR3;
  logic [31:0] zll_quarterround_quarterround25_outR3;
  logic [63:0] binop_inR7;
  logic [127:0] zll_quarterround_quarterround30_in;
  assign zll_quarterround_quarterround34_in = arg0;
  assign zll_quarterround_quarterround2_in = {zll_quarterround_quarterround34_in[63:32], zll_quarterround_quarterround34_in[127:96], zll_quarterround_quarterround34_in[95:64], zll_quarterround_quarterround34_in[31:0]};
  assign binop_in = {zll_quarterround_quarterround2_in[95:64], zll_quarterround_quarterround2_in[31:0]};
  assign zll_quarterround_quarterround28_in = binop_in[63:32] + binop_in[31:0];
  assign zll_quarterround_quarterround25_in = {32'h7, zll_quarterround_quarterround28_in[31:0]};
  ZLL_QuarterRound_quarterround25  inst (zll_quarterround_quarterround25_in[63:0], zll_quarterround_quarterround25_out);
  assign binop_inR1 = {zll_quarterround_quarterround2_in[63:32], zll_quarterround_quarterround25_out};
  assign zll_quarterround_quarterround16_in = {zll_quarterround_quarterround2_in[127:96], zll_quarterround_quarterround2_in[95:64], zll_quarterround_quarterround2_in[31:0], binop_inR1[63:32] ^ binop_inR1[31:0]};
  assign binop_inR2 = {zll_quarterround_quarterround16_in[31:0], zll_quarterround_quarterround16_in[95:64]};
  assign zll_quarterround_quarterround4_in = binop_inR2[63:32] + binop_inR2[31:0];
  assign zll_quarterround_quarterround25_inR1 = {32'h9, zll_quarterround_quarterround4_in[31:0]};
  ZLL_QuarterRound_quarterround25  instR1 (zll_quarterround_quarterround25_inR1[63:0], zll_quarterround_quarterround25_outR1);
  assign binop_inR3 = {zll_quarterround_quarterround16_in[127:96], zll_quarterround_quarterround25_outR1};
  assign zll_quarterround_quarterround40_in = {zll_quarterround_quarterround16_in[95:64], zll_quarterround_quarterround16_in[31:0], zll_quarterround_quarterround16_in[63:32], binop_inR3[63:32] ^ binop_inR3[31:0]};
  assign binop_inR4 = {zll_quarterround_quarterround40_in[31:0], zll_quarterround_quarterround40_in[95:64]};
  assign zll_quarterround_quarterround12_in = binop_inR4[63:32] + binop_inR4[31:0];
  assign zll_quarterround_quarterround25_inR2 = {32'hd, zll_quarterround_quarterround12_in[31:0]};
  ZLL_QuarterRound_quarterround25  instR2 (zll_quarterround_quarterround25_inR2[63:0], zll_quarterround_quarterround25_outR2);
  assign binop_inR5 = {zll_quarterround_quarterround40_in[63:32], zll_quarterround_quarterround25_outR2};
  assign zll_quarterround_quarterround6_in = {zll_quarterround_quarterround40_in[31:0], zll_quarterround_quarterround40_in[127:96], zll_quarterround_quarterround40_in[95:64], binop_inR5[63:32] ^ binop_inR5[31:0]};
  assign binop_inR6 = {zll_quarterround_quarterround6_in[31:0], zll_quarterround_quarterround6_in[127:96]};
  assign zll_quarterround_quarterround17_in = binop_inR6[63:32] + binop_inR6[31:0];
  assign zll_quarterround_quarterround25_inR3 = {32'h12, zll_quarterround_quarterround17_in[31:0]};
  ZLL_QuarterRound_quarterround25  instR3 (zll_quarterround_quarterround25_inR3[63:0], zll_quarterround_quarterround25_outR3);
  assign binop_inR7 = {zll_quarterround_quarterround6_in[95:64], zll_quarterround_quarterround25_outR3};
  assign zll_quarterround_quarterround30_in = {zll_quarterround_quarterround6_in[127:96], zll_quarterround_quarterround6_in[63:32], zll_quarterround_quarterround6_in[31:0], binop_inR7[63:32] ^ binop_inR7[31:0]};
  assign res = {zll_quarterround_quarterround30_in[31:0], zll_quarterround_quarterround30_in[95:64], zll_quarterround_quarterround30_in[127:96], zll_quarterround_quarterround30_in[63:32]};
endmodule

module Main_refold2 (input logic [5129:0] arg0,
  input logic [512:0] arg1,
  output logic [6157:0] res);
  logic [5642:0] main_conn10_in;
  logic [5129:0] main_conn10_out;
  logic [5129:0] zll_main_ten11_in;
  logic [5129:0] zll_main_ten11_out;
  logic [5129:0] zll_main_out101_in;
  logic [512:0] zll_main_out101_out;
  assign main_conn10_in = {arg0, arg1};
  Main_conn10  inst (main_conn10_in[5642:513], main_conn10_in[512:0], main_conn10_out);
  assign zll_main_ten11_in = main_conn10_out;
  ZLL_Main_ten11  instR1 (zll_main_ten11_in[5129:0], zll_main_ten11_out);
  assign zll_main_out101_in = zll_main_ten11_out;
  ZLL_Main_out101  instR2 (zll_main_out101_in[5129:0], zll_main_out101_out);
  assign res = {zll_main_out101_out, 2'h0, arg1, arg0};
endmodule

module ZLL_Main_ten11 (input logic [5129:0] arg0,
  output logic [5129:0] res);
  logic [5129:0] zll_main_ten9_in;
  logic [5129:0] zll_main_ten4_in;
  logic [5129:0] zll_main_ten_in;
  logic [5129:0] zll_main_ten7_in;
  logic [5129:0] zll_main_ten10_in;
  logic [5129:0] zll_main_ten2_in;
  logic [5129:0] zll_main_ten5_in;
  logic [512:0] main_dr1_in;
  logic [512:0] main_dr1_out;
  logic [512:0] main_dr1_inR1;
  logic [512:0] main_dr1_outR1;
  logic [512:0] main_dr1_inR2;
  logic [512:0] main_dr1_outR2;
  logic [512:0] main_dr1_inR3;
  logic [512:0] main_dr1_outR3;
  logic [512:0] main_dr1_inR4;
  logic [512:0] main_dr1_outR4;
  logic [512:0] main_dr1_inR5;
  logic [512:0] main_dr1_outR5;
  logic [512:0] main_dr1_inR6;
  logic [512:0] main_dr1_outR6;
  logic [512:0] main_dr1_inR7;
  logic [512:0] main_dr1_outR7;
  logic [512:0] main_dr1_inR8;
  logic [512:0] main_dr1_outR8;
  logic [512:0] main_dr1_inR9;
  logic [512:0] main_dr1_outR9;
  assign zll_main_ten9_in = arg0;
  assign zll_main_ten4_in = {zll_main_ten9_in[5129:4617], zll_main_ten9_in[3590:3078], zll_main_ten9_in[4616:4104], zll_main_ten9_in[4103:3591], zll_main_ten9_in[3077:2565], zll_main_ten9_in[2564:2052], zll_main_ten9_in[2051:1539], zll_main_ten9_in[1538:1026], zll_main_ten9_in[1025:513], zll_main_ten9_in[512:0]};
  assign zll_main_ten_in = {zll_main_ten4_in[3077:2565], zll_main_ten4_in[5129:4617], zll_main_ten4_in[4616:4104], zll_main_ten4_in[4103:3591], zll_main_ten4_in[3590:3078], zll_main_ten4_in[2564:2052], zll_main_ten4_in[2051:1539], zll_main_ten4_in[1538:1026], zll_main_ten4_in[1025:513], zll_main_ten4_in[512:0]};
  assign zll_main_ten7_in = {zll_main_ten_in[5129:4617], zll_main_ten_in[4616:4104], zll_main_ten_in[4103:3591], zll_main_ten_in[2564:2052], zll_main_ten_in[3590:3078], zll_main_ten_in[3077:2565], zll_main_ten_in[2051:1539], zll_main_ten_in[1538:1026], zll_main_ten_in[1025:513], zll_main_ten_in[512:0]};
  assign zll_main_ten10_in = {zll_main_ten7_in[5129:4617], zll_main_ten7_in[4616:4104], zll_main_ten7_in[2051:1539], zll_main_ten7_in[4103:3591], zll_main_ten7_in[3590:3078], zll_main_ten7_in[3077:2565], zll_main_ten7_in[2564:2052], zll_main_ten7_in[1538:1026], zll_main_ten7_in[1025:513], zll_main_ten7_in[512:0]};
  assign zll_main_ten2_in = {zll_main_ten10_in[5129:4617], zll_main_ten10_in[4616:4104], zll_main_ten10_in[4103:3591], zll_main_ten10_in[1538:1026], zll_main_ten10_in[3590:3078], zll_main_ten10_in[3077:2565], zll_main_ten10_in[2564:2052], zll_main_ten10_in[2051:1539], zll_main_ten10_in[1025:513], zll_main_ten10_in[512:0]};
  assign zll_main_ten5_in = {zll_main_ten2_in[5129:4617], zll_main_ten2_in[1025:513], zll_main_ten2_in[4616:4104], zll_main_ten2_in[4103:3591], zll_main_ten2_in[3590:3078], zll_main_ten2_in[3077:2565], zll_main_ten2_in[2564:2052], zll_main_ten2_in[2051:1539], zll_main_ten2_in[1538:1026], zll_main_ten2_in[512:0]};
  assign main_dr1_in = zll_main_ten5_in[4103:3591];
  Main_dr1  inst (main_dr1_in[512:0], main_dr1_out);
  assign main_dr1_inR1 = zll_main_ten5_in[1538:1026];
  Main_dr1  instR1 (main_dr1_inR1[512:0], main_dr1_outR1);
  assign main_dr1_inR2 = zll_main_ten5_in[1025:513];
  Main_dr1  instR2 (main_dr1_inR2[512:0], main_dr1_outR2);
  assign main_dr1_inR3 = zll_main_ten5_in[2564:2052];
  Main_dr1  instR3 (main_dr1_inR3[512:0], main_dr1_outR3);
  assign main_dr1_inR4 = zll_main_ten5_in[5129:4617];
  Main_dr1  instR4 (main_dr1_inR4[512:0], main_dr1_outR4);
  assign main_dr1_inR5 = zll_main_ten5_in[2051:1539];
  Main_dr1  instR5 (main_dr1_inR5[512:0], main_dr1_outR5);
  assign main_dr1_inR6 = zll_main_ten5_in[3590:3078];
  Main_dr1  instR6 (main_dr1_inR6[512:0], main_dr1_outR6);
  assign main_dr1_inR7 = zll_main_ten5_in[3077:2565];
  Main_dr1  instR7 (main_dr1_inR7[512:0], main_dr1_outR7);
  assign main_dr1_inR8 = zll_main_ten5_in[4616:4104];
  Main_dr1  instR8 (main_dr1_inR8[512:0], main_dr1_outR8);
  assign main_dr1_inR9 = zll_main_ten5_in[512:0];
  Main_dr1  instR9 (main_dr1_inR9[512:0], main_dr1_outR9);
  assign res = {main_dr1_out, main_dr1_outR1, main_dr1_outR2, main_dr1_outR3, main_dr1_outR4, main_dr1_outR5, main_dr1_outR6, main_dr1_outR7, main_dr1_outR8, main_dr1_outR9};
endmodule

module ZLL_QuarterRound_quarterround25 (input logic [63:0] arg0,
  output logic [31:0] res);
  logic [63:0] zll_quarterround_quarterround41_in;
  logic [63:0] binop_in;
  logic [63:0] binop_inR1;
  logic [63:0] binop_inR2;
  logic [63:0] binop_inR3;
  assign zll_quarterround_quarterround41_in = arg0;
  assign binop_in = {zll_quarterround_quarterround41_in[31:0], zll_quarterround_quarterround41_in[63:32]};
  assign binop_inR1 = {32'h20, zll_quarterround_quarterround41_in[63:32]};
  assign binop_inR2 = {zll_quarterround_quarterround41_in[31:0], binop_inR1[63:32] - binop_inR1[31:0]};
  assign binop_inR3 = {binop_in[63:32] << binop_in[31:0], binop_inR2[63:32] >> binop_inR2[31:0]};
  assign res = binop_inR3[63:32] | binop_inR3[31:0];
endmodule

module Main_dr1 (input logic [512:0] arg0,
  output logic [512:0] res);
  logic [1025:0] zll_main_dr12_in;
  logic [512:0] zll_main_dr1_in;
  logic [512:0] zll_main_dr11_in;
  logic [511:0] zll_columnround_columnround6_in;
  logic [511:0] zll_columnround_columnround11_in;
  logic [511:0] zll_columnround_columnround_in;
  logic [511:0] zll_columnround_columnround25_in;
  logic [511:0] zll_columnround_columnround21_in;
  logic [511:0] zll_columnround_columnround14_in;
  logic [511:0] zll_columnround_columnround16_in;
  logic [511:0] zll_columnround_columnround4_in;
  logic [511:0] zll_columnround_columnround28_in;
  logic [511:0] zll_columnround_columnround23_in;
  logic [511:0] zll_columnround_columnround29_in;
  logic [511:0] zll_columnround_columnround33_in;
  logic [511:0] zll_columnround_columnround17_in;
  logic [511:0] zll_columnround_columnround37_in;
  logic [511:0] zll_columnround_columnround9_in;
  logic [127:0] zll_quarterround_quarterround39_in;
  logic [127:0] zll_quarterround_quarterround39_out;
  logic [511:0] zll_columnround_columnround13_in;
  logic [511:0] zll_columnround_columnround32_in;
  logic [511:0] zll_columnround_columnround12_in;
  logic [511:0] zll_columnround_columnround2_in;
  logic [511:0] zll_columnround_columnround10_in;
  logic [127:0] zll_quarterround_quarterround39_inR1;
  logic [127:0] zll_quarterround_quarterround39_outR1;
  logic [511:0] zll_columnround_columnround8_in;
  logic [511:0] zll_columnround_columnround31_in;
  logic [511:0] zll_columnround_columnround5_in;
  logic [511:0] zll_columnround_columnround20_in;
  logic [127:0] zll_quarterround_quarterround39_inR2;
  logic [127:0] zll_quarterround_quarterround39_outR2;
  logic [511:0] zll_columnround_columnround30_in;
  logic [511:0] zll_columnround_columnround38_in;
  logic [511:0] zll_columnround_columnround22_in;
  logic [511:0] zll_columnround_columnround18_in;
  logic [511:0] zll_columnround_columnround34_in;
  logic [127:0] zll_quarterround_quarterround39_inR3;
  logic [127:0] zll_quarterround_quarterround39_outR3;
  logic [511:0] zll_columnround_columnround36_in;
  logic [511:0] zll_columnround_columnround19_in;
  logic [511:0] zll_columnround_columnround35_in;
  logic [511:0] zll_columnround_columnround3_in;
  logic [511:0] zll_columnround_columnround27_in;
  logic [511:0] zll_rowround_rowround36_in;
  logic [511:0] zll_rowround_rowround4_in;
  logic [511:0] zll_rowround_rowround20_in;
  logic [511:0] zll_rowround_rowround16_in;
  logic [511:0] zll_rowround_rowround24_in;
  logic [511:0] zll_rowround_rowround18_in;
  logic [511:0] zll_rowround_rowround37_in;
  logic [511:0] zll_rowround_rowround29_in;
  logic [511:0] zll_rowround_rowround9_in;
  logic [511:0] zll_rowround_rowround28_in;
  logic [511:0] zll_rowround_rowround35_in;
  logic [511:0] zll_rowround_rowround26_in;
  logic [511:0] zll_rowround_rowround19_in;
  logic [511:0] zll_rowround_rowround6_in;
  logic [127:0] zll_quarterround_quarterround39_inR4;
  logic [127:0] zll_quarterround_quarterround39_outR4;
  logic [511:0] zll_rowround_rowround17_in;
  logic [511:0] zll_rowround_rowround32_in;
  logic [511:0] zll_rowround_rowround31_in;
  logic [511:0] zll_rowround_rowround33_in;
  logic [127:0] zll_quarterround_quarterround39_inR5;
  logic [127:0] zll_quarterround_quarterround39_outR5;
  logic [511:0] zll_rowround_rowround25_in;
  logic [511:0] zll_rowround_rowround14_in;
  logic [511:0] zll_rowround_rowround7_in;
  logic [511:0] zll_rowround_rowround13_in;
  logic [511:0] zll_rowround_rowround11_in;
  logic [127:0] zll_quarterround_quarterround39_inR6;
  logic [127:0] zll_quarterround_quarterround39_outR6;
  logic [511:0] zll_rowround_rowround2_in;
  logic [511:0] zll_rowround_rowround8_in;
  logic [511:0] zll_rowround_rowround12_in;
  logic [511:0] zll_rowround_rowround5_in;
  logic [511:0] zll_rowround_rowround1_in;
  logic [127:0] zll_quarterround_quarterround39_inR7;
  logic [127:0] zll_quarterround_quarterround39_outR7;
  logic [511:0] zll_rowround_rowround21_in;
  logic [511:0] zll_rowround_rowround39_in;
  logic [511:0] zll_rowround_rowround27_in;
  logic [511:0] zll_rowround_rowround10_in;
  logic [512:0] lit_in;
  assign zll_main_dr12_in = {arg0, arg0};
  assign zll_main_dr1_in = zll_main_dr12_in[1025:513];
  assign zll_main_dr11_in = zll_main_dr1_in[512:0];
  assign zll_columnround_columnround6_in = zll_main_dr11_in[511:0];
  assign zll_columnround_columnround11_in = zll_columnround_columnround6_in[511:0];
  assign zll_columnround_columnround_in = {zll_columnround_columnround11_in[511:480], zll_columnround_columnround11_in[447:416], zll_columnround_columnround11_in[479:448], zll_columnround_columnround11_in[415:384], zll_columnround_columnround11_in[383:352], zll_columnround_columnround11_in[351:320], zll_columnround_columnround11_in[319:288], zll_columnround_columnround11_in[287:256], zll_columnround_columnround11_in[255:224], zll_columnround_columnround11_in[223:192], zll_columnround_columnround11_in[191:160], zll_columnround_columnround11_in[159:128], zll_columnround_columnround11_in[127:96], zll_columnround_columnround11_in[95:64], zll_columnround_columnround11_in[63:32], zll_columnround_columnround11_in[31:0]};
  assign zll_columnround_columnround25_in = {zll_columnround_columnround_in[511:480], zll_columnround_columnround_in[415:384], zll_columnround_columnround_in[479:448], zll_columnround_columnround_in[447:416], zll_columnround_columnround_in[383:352], zll_columnround_columnround_in[351:320], zll_columnround_columnround_in[319:288], zll_columnround_columnround_in[287:256], zll_columnround_columnround_in[255:224], zll_columnround_columnround_in[223:192], zll_columnround_columnround_in[191:160], zll_columnround_columnround_in[159:128], zll_columnround_columnround_in[127:96], zll_columnround_columnround_in[95:64], zll_columnround_columnround_in[63:32], zll_columnround_columnround_in[31:0]};
  assign zll_columnround_columnround21_in = {zll_columnround_columnround25_in[511:480], zll_columnround_columnround25_in[383:352], zll_columnround_columnround25_in[479:448], zll_columnround_columnround25_in[447:416], zll_columnround_columnround25_in[415:384], zll_columnround_columnround25_in[351:320], zll_columnround_columnround25_in[319:288], zll_columnround_columnround25_in[287:256], zll_columnround_columnround25_in[255:224], zll_columnround_columnround25_in[223:192], zll_columnround_columnround25_in[191:160], zll_columnround_columnround25_in[159:128], zll_columnround_columnround25_in[127:96], zll_columnround_columnround25_in[95:64], zll_columnround_columnround25_in[63:32], zll_columnround_columnround25_in[31:0]};
  assign zll_columnround_columnround14_in = {zll_columnround_columnround21_in[511:480], zll_columnround_columnround21_in[351:320], zll_columnround_columnround21_in[479:448], zll_columnround_columnround21_in[447:416], zll_columnround_columnround21_in[415:384], zll_columnround_columnround21_in[383:352], zll_columnround_columnround21_in[319:288], zll_columnround_columnround21_in[287:256], zll_columnround_columnround21_in[255:224], zll_columnround_columnround21_in[223:192], zll_columnround_columnround21_in[191:160], zll_columnround_columnround21_in[159:128], zll_columnround_columnround21_in[127:96], zll_columnround_columnround21_in[95:64], zll_columnround_columnround21_in[63:32], zll_columnround_columnround21_in[31:0]};
  assign zll_columnround_columnround16_in = {zll_columnround_columnround14_in[319:288], zll_columnround_columnround14_in[511:480], zll_columnround_columnround14_in[479:448], zll_columnround_columnround14_in[447:416], zll_columnround_columnround14_in[415:384], zll_columnround_columnround14_in[383:352], zll_columnround_columnround14_in[351:320], zll_columnround_columnround14_in[287:256], zll_columnround_columnround14_in[255:224], zll_columnround_columnround14_in[223:192], zll_columnround_columnround14_in[191:160], zll_columnround_columnround14_in[159:128], zll_columnround_columnround14_in[127:96], zll_columnround_columnround14_in[95:64], zll_columnround_columnround14_in[63:32], zll_columnround_columnround14_in[31:0]};
  assign zll_columnround_columnround4_in = {zll_columnround_columnround16_in[511:480], zll_columnround_columnround16_in[479:448], zll_columnround_columnround16_in[287:256], zll_columnround_columnround16_in[447:416], zll_columnround_columnround16_in[415:384], zll_columnround_columnround16_in[383:352], zll_columnround_columnround16_in[351:320], zll_columnround_columnround16_in[319:288], zll_columnround_columnround16_in[255:224], zll_columnround_columnround16_in[223:192], zll_columnround_columnround16_in[191:160], zll_columnround_columnround16_in[159:128], zll_columnround_columnround16_in[127:96], zll_columnround_columnround16_in[95:64], zll_columnround_columnround16_in[63:32], zll_columnround_columnround16_in[31:0]};
  assign zll_columnround_columnround28_in = {zll_columnround_columnround4_in[511:480], zll_columnround_columnround4_in[479:448], zll_columnround_columnround4_in[447:416], zll_columnround_columnround4_in[415:384], zll_columnround_columnround4_in[383:352], zll_columnround_columnround4_in[351:320], zll_columnround_columnround4_in[255:224], zll_columnround_columnround4_in[319:288], zll_columnround_columnround4_in[287:256], zll_columnround_columnround4_in[223:192], zll_columnround_columnround4_in[191:160], zll_columnround_columnround4_in[159:128], zll_columnround_columnround4_in[127:96], zll_columnround_columnround4_in[95:64], zll_columnround_columnround4_in[63:32], zll_columnround_columnround4_in[31:0]};
  assign zll_columnround_columnround23_in = {zll_columnround_columnround28_in[511:480], zll_columnround_columnround28_in[223:192], zll_columnround_columnround28_in[479:448], zll_columnround_columnround28_in[447:416], zll_columnround_columnround28_in[415:384], zll_columnround_columnround28_in[383:352], zll_columnround_columnround28_in[351:320], zll_columnround_columnround28_in[319:288], zll_columnround_columnround28_in[287:256], zll_columnround_columnround28_in[255:224], zll_columnround_columnround28_in[191:160], zll_columnround_columnround28_in[159:128], zll_columnround_columnround28_in[127:96], zll_columnround_columnround28_in[95:64], zll_columnround_columnround28_in[63:32], zll_columnround_columnround28_in[31:0]};
  assign zll_columnround_columnround29_in = {zll_columnround_columnround23_in[511:480], zll_columnround_columnround23_in[191:160], zll_columnround_columnround23_in[479:448], zll_columnround_columnround23_in[447:416], zll_columnround_columnround23_in[415:384], zll_columnround_columnround23_in[383:352], zll_columnround_columnround23_in[351:320], zll_columnround_columnround23_in[319:288], zll_columnround_columnround23_in[287:256], zll_columnround_columnround23_in[255:224], zll_columnround_columnround23_in[223:192], zll_columnround_columnround23_in[159:128], zll_columnround_columnround23_in[127:96], zll_columnround_columnround23_in[95:64], zll_columnround_columnround23_in[63:32], zll_columnround_columnround23_in[31:0]};
  assign zll_columnround_columnround33_in = {zll_columnround_columnround29_in[511:480], zll_columnround_columnround29_in[479:448], zll_columnround_columnround29_in[159:128], zll_columnround_columnround29_in[447:416], zll_columnround_columnround29_in[415:384], zll_columnround_columnround29_in[383:352], zll_columnround_columnround29_in[351:320], zll_columnround_columnround29_in[319:288], zll_columnround_columnround29_in[287:256], zll_columnround_columnround29_in[255:224], zll_columnround_columnround29_in[223:192], zll_columnround_columnround29_in[191:160], zll_columnround_columnround29_in[127:96], zll_columnround_columnround29_in[95:64], zll_columnround_columnround29_in[63:32], zll_columnround_columnround29_in[31:0]};
  assign zll_columnround_columnround17_in = {zll_columnround_columnround33_in[511:480], zll_columnround_columnround33_in[127:96], zll_columnround_columnround33_in[479:448], zll_columnround_columnround33_in[447:416], zll_columnround_columnround33_in[415:384], zll_columnround_columnround33_in[383:352], zll_columnround_columnround33_in[351:320], zll_columnround_columnround33_in[319:288], zll_columnround_columnround33_in[287:256], zll_columnround_columnround33_in[255:224], zll_columnround_columnround33_in[223:192], zll_columnround_columnround33_in[191:160], zll_columnround_columnround33_in[159:128], zll_columnround_columnround33_in[95:64], zll_columnround_columnround33_in[63:32], zll_columnround_columnround33_in[31:0]};
  assign zll_columnround_columnround37_in = {zll_columnround_columnround17_in[511:480], zll_columnround_columnround17_in[479:448], zll_columnround_columnround17_in[447:416], zll_columnround_columnround17_in[415:384], zll_columnround_columnround17_in[383:352], zll_columnround_columnround17_in[351:320], zll_columnround_columnround17_in[319:288], zll_columnround_columnround17_in[287:256], zll_columnround_columnround17_in[255:224], zll_columnround_columnround17_in[95:64], zll_columnround_columnround17_in[223:192], zll_columnround_columnround17_in[191:160], zll_columnround_columnround17_in[159:128], zll_columnround_columnround17_in[127:96], zll_columnround_columnround17_in[63:32], zll_columnround_columnround17_in[31:0]};
  assign zll_columnround_columnround9_in = {zll_columnround_columnround37_in[511:480], zll_columnround_columnround37_in[479:448], zll_columnround_columnround37_in[447:416], zll_columnround_columnround37_in[63:32], zll_columnround_columnround37_in[415:384], zll_columnround_columnround37_in[383:352], zll_columnround_columnround37_in[351:320], zll_columnround_columnround37_in[319:288], zll_columnround_columnround37_in[287:256], zll_columnround_columnround37_in[255:224], zll_columnround_columnround37_in[223:192], zll_columnround_columnround37_in[191:160], zll_columnround_columnround37_in[159:128], zll_columnround_columnround37_in[127:96], zll_columnround_columnround37_in[95:64], zll_columnround_columnround37_in[31:0]};
  assign zll_quarterround_quarterround39_in = {zll_columnround_columnround9_in[319:288], zll_columnround_columnround9_in[223:192], zll_columnround_columnround9_in[127:96], zll_columnround_columnround9_in[479:448]};
  ZLL_QuarterRound_quarterround39  inst (zll_quarterround_quarterround39_in[127:0], zll_quarterround_quarterround39_out);
  assign zll_columnround_columnround13_in = {zll_columnround_columnround9_in[511:480], zll_columnround_columnround9_in[31:0], zll_columnround_columnround9_in[447:416], zll_columnround_columnround9_in[415:384], zll_columnround_columnround9_in[383:352], zll_columnround_columnround9_in[351:320], zll_columnround_columnround9_in[287:256], zll_columnround_columnround9_in[255:224], zll_columnround_columnround9_in[191:160], zll_columnround_columnround9_in[159:128], zll_columnround_columnround9_in[95:64], zll_columnround_columnround9_in[63:32], zll_quarterround_quarterround39_out};
  assign zll_columnround_columnround32_in = {zll_columnround_columnround13_in[511:480], zll_columnround_columnround13_in[479:448], zll_columnround_columnround13_in[447:416], zll_columnround_columnround13_in[415:384], zll_columnround_columnround13_in[383:352], zll_columnround_columnround13_in[351:320], zll_columnround_columnround13_in[319:288], zll_columnround_columnround13_in[287:256], zll_columnround_columnround13_in[255:224], zll_columnround_columnround13_in[223:192], zll_columnround_columnround13_in[191:160], zll_columnround_columnround13_in[159:128], zll_columnround_columnround13_in[127:0]};
  assign zll_columnround_columnround12_in = {zll_columnround_columnround32_in[511:480], zll_columnround_columnround32_in[127:96], zll_columnround_columnround32_in[479:448], zll_columnround_columnround32_in[447:416], zll_columnround_columnround32_in[415:384], zll_columnround_columnround32_in[383:352], zll_columnround_columnround32_in[351:320], zll_columnround_columnround32_in[319:288], zll_columnround_columnround32_in[287:256], zll_columnround_columnround32_in[255:224], zll_columnround_columnround32_in[223:192], zll_columnround_columnround32_in[191:160], zll_columnround_columnround32_in[159:128], zll_columnround_columnround32_in[95:64], zll_columnround_columnround32_in[63:32], zll_columnround_columnround32_in[31:0]};
  assign zll_columnround_columnround2_in = {zll_columnround_columnround12_in[511:480], zll_columnround_columnround12_in[479:448], zll_columnround_columnround12_in[447:416], zll_columnround_columnround12_in[415:384], zll_columnround_columnround12_in[383:352], zll_columnround_columnround12_in[351:320], zll_columnround_columnround12_in[319:288], zll_columnround_columnround12_in[287:256], zll_columnround_columnround12_in[255:224], zll_columnround_columnround12_in[223:192], zll_columnround_columnround12_in[191:160], zll_columnround_columnround12_in[95:64], zll_columnround_columnround12_in[159:128], zll_columnround_columnround12_in[127:96], zll_columnround_columnround12_in[63:32], zll_columnround_columnround12_in[31:0]};
  assign zll_columnround_columnround10_in = {zll_columnround_columnround2_in[511:480], zll_columnround_columnround2_in[479:448], zll_columnround_columnround2_in[447:416], zll_columnround_columnround2_in[415:384], zll_columnround_columnround2_in[383:352], zll_columnround_columnround2_in[351:320], zll_columnround_columnround2_in[319:288], zll_columnround_columnround2_in[63:32], zll_columnround_columnround2_in[287:256], zll_columnround_columnround2_in[255:224], zll_columnround_columnround2_in[223:192], zll_columnround_columnround2_in[191:160], zll_columnround_columnround2_in[159:128], zll_columnround_columnround2_in[127:96], zll_columnround_columnround2_in[95:64], zll_columnround_columnround2_in[31:0]};
  assign zll_quarterround_quarterround39_inR1 = {zll_columnround_columnround10_in[223:192], zll_columnround_columnround10_in[319:288], zll_columnround_columnround10_in[191:160], zll_columnround_columnround10_in[63:32]};
  ZLL_QuarterRound_quarterround39  instR1 (zll_quarterround_quarterround39_inR1[127:0], zll_quarterround_quarterround39_outR1);
  assign zll_columnround_columnround8_in = {zll_columnround_columnround10_in[511:480], zll_columnround_columnround10_in[31:0], zll_columnround_columnround10_in[479:448], zll_columnround_columnround10_in[447:416], zll_columnround_columnround10_in[415:384], zll_columnround_columnround10_in[383:352], zll_columnround_columnround10_in[351:320], zll_columnround_columnround10_in[287:256], zll_columnround_columnround10_in[255:224], zll_columnround_columnround10_in[159:128], zll_columnround_columnround10_in[127:96], zll_columnround_columnround10_in[95:64], zll_quarterround_quarterround39_outR1};
  assign zll_columnround_columnround31_in = {zll_columnround_columnround8_in[511:480], zll_columnround_columnround8_in[479:448], zll_columnround_columnround8_in[447:416], zll_columnround_columnround8_in[415:384], zll_columnround_columnround8_in[383:352], zll_columnround_columnround8_in[351:320], zll_columnround_columnround8_in[319:288], zll_columnround_columnround8_in[287:256], zll_columnround_columnround8_in[255:224], zll_columnround_columnround8_in[223:192], zll_columnround_columnround8_in[191:160], zll_columnround_columnround8_in[159:128], zll_columnround_columnround8_in[127:0]};
  assign zll_columnround_columnround5_in = {zll_columnround_columnround31_in[511:480], zll_columnround_columnround31_in[479:448], zll_columnround_columnround31_in[447:416], zll_columnround_columnround31_in[415:384], zll_columnround_columnround31_in[383:352], zll_columnround_columnround31_in[351:320], zll_columnround_columnround31_in[319:288], zll_columnround_columnround31_in[127:96], zll_columnround_columnround31_in[287:256], zll_columnround_columnround31_in[255:224], zll_columnround_columnround31_in[223:192], zll_columnround_columnround31_in[191:160], zll_columnround_columnround31_in[159:128], zll_columnround_columnround31_in[95:64], zll_columnround_columnround31_in[63:32], zll_columnround_columnround31_in[31:0]};
  assign zll_columnround_columnround20_in = {zll_columnround_columnround5_in[511:480], zll_columnround_columnround5_in[479:448], zll_columnround_columnround5_in[447:416], zll_columnround_columnround5_in[415:384], zll_columnround_columnround5_in[383:352], zll_columnround_columnround5_in[351:320], zll_columnround_columnround5_in[319:288], zll_columnround_columnround5_in[287:256], zll_columnround_columnround5_in[255:224], zll_columnround_columnround5_in[223:192], zll_columnround_columnround5_in[63:32], zll_columnround_columnround5_in[191:160], zll_columnround_columnround5_in[159:128], zll_columnround_columnround5_in[127:96], zll_columnround_columnround5_in[95:64], zll_columnround_columnround5_in[31:0]};
  assign zll_quarterround_quarterround39_inR2 = {zll_columnround_columnround20_in[383:352], zll_columnround_columnround20_in[351:320], zll_columnround_columnround20_in[95:64], zll_columnround_columnround20_in[511:480]};
  ZLL_QuarterRound_quarterround39  instR2 (zll_quarterround_quarterround39_inR2[127:0], zll_quarterround_quarterround39_outR2);
  assign zll_columnround_columnround30_in = {zll_columnround_columnround20_in[479:448], zll_columnround_columnround20_in[447:416], zll_columnround_columnround20_in[415:384], zll_columnround_columnround20_in[319:288], zll_columnround_columnround20_in[287:256], zll_columnround_columnround20_in[255:224], zll_columnround_columnround20_in[223:192], zll_columnround_columnround20_in[31:0], zll_columnround_columnround20_in[191:160], zll_columnround_columnround20_in[159:128], zll_columnround_columnround20_in[127:96], zll_columnround_columnround20_in[63:32], zll_quarterround_quarterround39_outR2};
  assign zll_columnround_columnround38_in = {zll_columnround_columnround30_in[511:480], zll_columnround_columnround30_in[479:448], zll_columnround_columnround30_in[447:416], zll_columnround_columnround30_in[415:384], zll_columnround_columnround30_in[383:352], zll_columnround_columnround30_in[351:320], zll_columnround_columnround30_in[319:288], zll_columnround_columnround30_in[287:256], zll_columnround_columnround30_in[255:224], zll_columnround_columnround30_in[223:192], zll_columnround_columnround30_in[191:160], zll_columnround_columnround30_in[159:128], zll_columnround_columnround30_in[127:0]};
  assign zll_columnround_columnround22_in = {zll_columnround_columnround38_in[511:480], zll_columnround_columnround38_in[479:448], zll_columnround_columnround38_in[447:416], zll_columnround_columnround38_in[415:384], zll_columnround_columnround38_in[383:352], zll_columnround_columnround38_in[351:320], zll_columnround_columnround38_in[319:288], zll_columnround_columnround38_in[287:256], zll_columnround_columnround38_in[255:224], zll_columnround_columnround38_in[223:192], zll_columnround_columnround38_in[127:96], zll_columnround_columnround38_in[191:160], zll_columnround_columnround38_in[159:128], zll_columnround_columnround38_in[95:64], zll_columnround_columnround38_in[63:32], zll_columnround_columnround38_in[31:0]};
  assign zll_columnround_columnround18_in = {zll_columnround_columnround22_in[511:480], zll_columnround_columnround22_in[479:448], zll_columnround_columnround22_in[447:416], zll_columnround_columnround22_in[415:384], zll_columnround_columnround22_in[383:352], zll_columnround_columnround22_in[351:320], zll_columnround_columnround22_in[319:288], zll_columnround_columnround22_in[287:256], zll_columnround_columnround22_in[255:224], zll_columnround_columnround22_in[223:192], zll_columnround_columnround22_in[191:160], zll_columnround_columnround22_in[159:128], zll_columnround_columnround22_in[95:64], zll_columnround_columnround22_in[127:96], zll_columnround_columnround22_in[63:32], zll_columnround_columnround22_in[31:0]};
  assign zll_columnround_columnround34_in = {zll_columnround_columnround18_in[511:480], zll_columnround_columnround18_in[479:448], zll_columnround_columnround18_in[447:416], zll_columnround_columnround18_in[415:384], zll_columnround_columnround18_in[383:352], zll_columnround_columnround18_in[351:320], zll_columnround_columnround18_in[63:32], zll_columnround_columnround18_in[319:288], zll_columnround_columnround18_in[287:256], zll_columnround_columnround18_in[255:224], zll_columnround_columnround18_in[223:192], zll_columnround_columnround18_in[191:160], zll_columnround_columnround18_in[159:128], zll_columnround_columnround18_in[127:96], zll_columnround_columnround18_in[95:64], zll_columnround_columnround18_in[31:0]};
  assign zll_quarterround_quarterround39_inR3 = {zll_columnround_columnround34_in[447:416], zll_columnround_columnround34_in[191:160], zll_columnround_columnround34_in[287:256], zll_columnround_columnround34_in[415:384]};
  ZLL_QuarterRound_quarterround39  instR3 (zll_quarterround_quarterround39_inR3[127:0], zll_quarterround_quarterround39_outR3);
  assign zll_columnround_columnround36_in = {zll_columnround_columnround34_in[511:480], zll_columnround_columnround34_in[31:0], zll_columnround_columnround34_in[479:448], zll_columnround_columnround34_in[383:352], zll_columnround_columnround34_in[351:320], zll_columnround_columnround34_in[319:288], zll_columnround_columnround34_in[255:224], zll_columnround_columnround34_in[223:192], zll_columnround_columnround34_in[159:128], zll_columnround_columnround34_in[127:96], zll_columnround_columnround34_in[95:64], zll_columnround_columnround34_in[63:32], zll_quarterround_quarterround39_outR3};
  assign zll_columnround_columnround19_in = {zll_columnround_columnround36_in[511:480], zll_columnround_columnround36_in[479:448], zll_columnround_columnround36_in[447:416], zll_columnround_columnround36_in[415:384], zll_columnround_columnround36_in[383:352], zll_columnround_columnround36_in[351:320], zll_columnround_columnround36_in[319:288], zll_columnround_columnround36_in[287:256], zll_columnround_columnround36_in[255:224], zll_columnround_columnround36_in[223:192], zll_columnround_columnround36_in[191:160], zll_columnround_columnround36_in[159:128], zll_columnround_columnround36_in[127:0]};
  assign zll_columnround_columnround35_in = {zll_columnround_columnround19_in[511:480], zll_columnround_columnround19_in[479:448], zll_columnround_columnround19_in[127:96], zll_columnround_columnround19_in[447:416], zll_columnround_columnround19_in[415:384], zll_columnround_columnround19_in[383:352], zll_columnround_columnround19_in[351:320], zll_columnround_columnround19_in[319:288], zll_columnround_columnround19_in[287:256], zll_columnround_columnround19_in[255:224], zll_columnround_columnround19_in[223:192], zll_columnround_columnround19_in[191:160], zll_columnround_columnround19_in[159:128], zll_columnround_columnround19_in[95:64], zll_columnround_columnround19_in[63:32], zll_columnround_columnround19_in[31:0]};
  assign zll_columnround_columnround3_in = {zll_columnround_columnround35_in[511:480], zll_columnround_columnround35_in[479:448], zll_columnround_columnround35_in[447:416], zll_columnround_columnround35_in[415:384], zll_columnround_columnround35_in[383:352], zll_columnround_columnround35_in[351:320], zll_columnround_columnround35_in[319:288], zll_columnround_columnround35_in[287:256], zll_columnround_columnround35_in[255:224], zll_columnround_columnround35_in[223:192], zll_columnround_columnround35_in[191:160], zll_columnround_columnround35_in[159:128], zll_columnround_columnround35_in[95:64], zll_columnround_columnround35_in[127:96], zll_columnround_columnround35_in[63:32], zll_columnround_columnround35_in[31:0]};
  assign zll_columnround_columnround27_in = {zll_columnround_columnround3_in[511:480], zll_columnround_columnround3_in[479:448], zll_columnround_columnround3_in[447:416], zll_columnround_columnround3_in[415:384], zll_columnround_columnround3_in[63:32], zll_columnround_columnround3_in[383:352], zll_columnround_columnround3_in[351:320], zll_columnround_columnround3_in[319:288], zll_columnround_columnround3_in[287:256], zll_columnround_columnround3_in[255:224], zll_columnround_columnround3_in[223:192], zll_columnround_columnround3_in[191:160], zll_columnround_columnround3_in[159:128], zll_columnround_columnround3_in[127:96], zll_columnround_columnround3_in[95:64], zll_columnround_columnround3_in[31:0]};
  assign zll_rowround_rowround36_in = {zll_columnround_columnround27_in[415:384], zll_columnround_columnround27_in[255:224], zll_columnround_columnround27_in[287:256], zll_columnround_columnround27_in[95:64], zll_columnround_columnround27_in[159:128], zll_columnround_columnround27_in[351:320], zll_columnround_columnround27_in[479:448], zll_columnround_columnround27_in[383:352], zll_columnround_columnround27_in[319:288], zll_columnround_columnround27_in[63:32], zll_columnround_columnround27_in[191:160], zll_columnround_columnround27_in[31:0], zll_columnround_columnround27_in[511:480], zll_columnround_columnround27_in[223:192], zll_columnround_columnround27_in[127:96], zll_columnround_columnround27_in[447:416]};
  assign zll_rowround_rowround4_in = zll_rowround_rowround36_in[511:0];
  assign zll_rowround_rowround20_in = {zll_rowround_rowround4_in[479:448], zll_rowround_rowround4_in[511:480], zll_rowround_rowround4_in[447:416], zll_rowround_rowround4_in[415:384], zll_rowround_rowround4_in[383:352], zll_rowround_rowround4_in[351:320], zll_rowround_rowround4_in[319:288], zll_rowround_rowround4_in[287:256], zll_rowround_rowround4_in[255:224], zll_rowround_rowround4_in[223:192], zll_rowround_rowround4_in[191:160], zll_rowround_rowround4_in[159:128], zll_rowround_rowround4_in[127:96], zll_rowround_rowround4_in[95:64], zll_rowround_rowround4_in[63:32], zll_rowround_rowround4_in[31:0]};
  assign zll_rowround_rowround16_in = {zll_rowround_rowround20_in[511:480], zll_rowround_rowround20_in[447:416], zll_rowround_rowround20_in[479:448], zll_rowround_rowround20_in[415:384], zll_rowround_rowround20_in[383:352], zll_rowround_rowround20_in[351:320], zll_rowround_rowround20_in[319:288], zll_rowround_rowround20_in[287:256], zll_rowround_rowround20_in[255:224], zll_rowround_rowround20_in[223:192], zll_rowround_rowround20_in[191:160], zll_rowround_rowround20_in[159:128], zll_rowround_rowround20_in[127:96], zll_rowround_rowround20_in[95:64], zll_rowround_rowround20_in[63:32], zll_rowround_rowround20_in[31:0]};
  assign zll_rowround_rowround24_in = {zll_rowround_rowround16_in[511:480], zll_rowround_rowround16_in[479:448], zll_rowround_rowround16_in[415:384], zll_rowround_rowround16_in[447:416], zll_rowround_rowround16_in[383:352], zll_rowround_rowround16_in[351:320], zll_rowround_rowround16_in[319:288], zll_rowround_rowround16_in[287:256], zll_rowround_rowround16_in[255:224], zll_rowround_rowround16_in[223:192], zll_rowround_rowround16_in[191:160], zll_rowround_rowround16_in[159:128], zll_rowround_rowround16_in[127:96], zll_rowround_rowround16_in[95:64], zll_rowround_rowround16_in[63:32], zll_rowround_rowround16_in[31:0]};
  assign zll_rowround_rowround18_in = {zll_rowround_rowround24_in[511:480], zll_rowround_rowround24_in[383:352], zll_rowround_rowround24_in[479:448], zll_rowround_rowround24_in[447:416], zll_rowround_rowround24_in[415:384], zll_rowround_rowround24_in[351:320], zll_rowround_rowround24_in[319:288], zll_rowround_rowround24_in[287:256], zll_rowround_rowround24_in[255:224], zll_rowround_rowround24_in[223:192], zll_rowround_rowround24_in[191:160], zll_rowround_rowround24_in[159:128], zll_rowround_rowround24_in[127:96], zll_rowround_rowround24_in[95:64], zll_rowround_rowround24_in[63:32], zll_rowround_rowround24_in[31:0]};
  assign zll_rowround_rowround37_in = {zll_rowround_rowround18_in[511:480], zll_rowround_rowround18_in[479:448], zll_rowround_rowround18_in[447:416], zll_rowround_rowround18_in[415:384], zll_rowround_rowround18_in[351:320], zll_rowround_rowround18_in[383:352], zll_rowround_rowround18_in[319:288], zll_rowround_rowround18_in[287:256], zll_rowround_rowround18_in[255:224], zll_rowround_rowround18_in[223:192], zll_rowround_rowround18_in[191:160], zll_rowround_rowround18_in[159:128], zll_rowround_rowround18_in[127:96], zll_rowround_rowround18_in[95:64], zll_rowround_rowround18_in[63:32], zll_rowround_rowround18_in[31:0]};
  assign zll_rowround_rowround29_in = {zll_rowround_rowround37_in[319:288], zll_rowround_rowround37_in[511:480], zll_rowround_rowround37_in[479:448], zll_rowround_rowround37_in[447:416], zll_rowround_rowround37_in[415:384], zll_rowround_rowround37_in[383:352], zll_rowround_rowround37_in[351:320], zll_rowround_rowround37_in[287:256], zll_rowround_rowround37_in[255:224], zll_rowround_rowround37_in[223:192], zll_rowround_rowround37_in[191:160], zll_rowround_rowround37_in[159:128], zll_rowround_rowround37_in[127:96], zll_rowround_rowround37_in[95:64], zll_rowround_rowround37_in[63:32], zll_rowround_rowround37_in[31:0]};
  assign zll_rowround_rowround9_in = {zll_rowround_rowround29_in[287:256], zll_rowround_rowround29_in[511:480], zll_rowround_rowround29_in[479:448], zll_rowround_rowround29_in[447:416], zll_rowround_rowround29_in[415:384], zll_rowround_rowround29_in[383:352], zll_rowround_rowround29_in[351:320], zll_rowround_rowround29_in[319:288], zll_rowround_rowround29_in[255:224], zll_rowround_rowround29_in[223:192], zll_rowround_rowround29_in[191:160], zll_rowround_rowround29_in[159:128], zll_rowround_rowround29_in[127:96], zll_rowround_rowround29_in[95:64], zll_rowround_rowround29_in[63:32], zll_rowround_rowround29_in[31:0]};
  assign zll_rowround_rowround28_in = {zll_rowround_rowround9_in[511:480], zll_rowround_rowround9_in[479:448], zll_rowround_rowround9_in[223:192], zll_rowround_rowround9_in[447:416], zll_rowround_rowround9_in[415:384], zll_rowround_rowround9_in[383:352], zll_rowround_rowround9_in[351:320], zll_rowround_rowround9_in[319:288], zll_rowround_rowround9_in[287:256], zll_rowround_rowround9_in[255:224], zll_rowround_rowround9_in[191:160], zll_rowround_rowround9_in[159:128], zll_rowround_rowround9_in[127:96], zll_rowround_rowround9_in[95:64], zll_rowround_rowround9_in[63:32], zll_rowround_rowround9_in[31:0]};
  assign zll_rowround_rowround35_in = {zll_rowround_rowround28_in[511:480], zll_rowround_rowround28_in[479:448], zll_rowround_rowround28_in[447:416], zll_rowround_rowround28_in[415:384], zll_rowround_rowround28_in[383:352], zll_rowround_rowround28_in[351:320], zll_rowround_rowround28_in[319:288], zll_rowround_rowround28_in[287:256], zll_rowround_rowround28_in[255:224], zll_rowround_rowround28_in[191:160], zll_rowround_rowround28_in[223:192], zll_rowround_rowround28_in[159:128], zll_rowround_rowround28_in[127:96], zll_rowround_rowround28_in[95:64], zll_rowround_rowround28_in[63:32], zll_rowround_rowround28_in[31:0]};
  assign zll_rowround_rowround26_in = {zll_rowround_rowround35_in[511:480], zll_rowround_rowround35_in[479:448], zll_rowround_rowround35_in[447:416], zll_rowround_rowround35_in[415:384], zll_rowround_rowround35_in[383:352], zll_rowround_rowround35_in[351:320], zll_rowround_rowround35_in[319:288], zll_rowround_rowround35_in[287:256], zll_rowround_rowround35_in[255:224], zll_rowround_rowround35_in[223:192], zll_rowround_rowround35_in[159:128], zll_rowround_rowround35_in[191:160], zll_rowround_rowround35_in[127:96], zll_rowround_rowround35_in[95:64], zll_rowround_rowround35_in[63:32], zll_rowround_rowround35_in[31:0]};
  assign zll_rowround_rowround19_in = {zll_rowround_rowround26_in[511:480], zll_rowround_rowround26_in[479:448], zll_rowround_rowround26_in[447:416], zll_rowround_rowround26_in[415:384], zll_rowround_rowround26_in[383:352], zll_rowround_rowround26_in[351:320], zll_rowround_rowround26_in[319:288], zll_rowround_rowround26_in[287:256], zll_rowround_rowround26_in[255:224], zll_rowround_rowround26_in[127:96], zll_rowround_rowround26_in[223:192], zll_rowround_rowround26_in[191:160], zll_rowround_rowround26_in[159:128], zll_rowround_rowround26_in[95:64], zll_rowround_rowround26_in[63:32], zll_rowround_rowround26_in[31:0]};
  assign zll_rowround_rowround6_in = {zll_rowround_rowround19_in[511:480], zll_rowround_rowround19_in[479:448], zll_rowround_rowround19_in[447:416], zll_rowround_rowround19_in[415:384], zll_rowround_rowround19_in[383:352], zll_rowround_rowround19_in[351:320], zll_rowround_rowround19_in[319:288], zll_rowround_rowround19_in[63:32], zll_rowround_rowround19_in[287:256], zll_rowround_rowround19_in[255:224], zll_rowround_rowround19_in[223:192], zll_rowround_rowround19_in[191:160], zll_rowround_rowround19_in[159:128], zll_rowround_rowround19_in[127:96], zll_rowround_rowround19_in[95:64], zll_rowround_rowround19_in[31:0]};
  assign zll_quarterround_quarterround39_inR4 = {zll_rowround_rowround6_in[223:192], zll_rowround_rowround6_in[415:384], zll_rowround_rowround6_in[351:320], zll_rowround_rowround6_in[319:288]};
  ZLL_QuarterRound_quarterround39  instR4 (zll_quarterround_quarterround39_inR4[127:0], zll_quarterround_quarterround39_outR4);
  assign zll_rowround_rowround17_in = {zll_rowround_rowround6_in[511:480], zll_rowround_rowround6_in[479:448], zll_rowround_rowround6_in[447:416], zll_rowround_rowround6_in[383:352], zll_rowround_rowround6_in[31:0], zll_rowround_rowround6_in[287:256], zll_rowround_rowround6_in[255:224], zll_rowround_rowround6_in[191:160], zll_rowround_rowround6_in[159:128], zll_rowround_rowround6_in[127:96], zll_rowround_rowround6_in[95:64], zll_rowround_rowround6_in[63:32], zll_quarterround_quarterround39_outR4};
  assign zll_rowround_rowround32_in = {zll_rowround_rowround17_in[511:480], zll_rowround_rowround17_in[479:448], zll_rowround_rowround17_in[447:416], zll_rowround_rowround17_in[415:384], zll_rowround_rowround17_in[383:352], zll_rowround_rowround17_in[351:320], zll_rowround_rowround17_in[319:288], zll_rowround_rowround17_in[287:256], zll_rowround_rowround17_in[255:224], zll_rowround_rowround17_in[223:192], zll_rowround_rowround17_in[191:160], zll_rowround_rowround17_in[159:128], zll_rowround_rowround17_in[127:0]};
  assign zll_rowround_rowround31_in = {zll_rowround_rowround32_in[511:480], zll_rowround_rowround32_in[479:448], zll_rowround_rowround32_in[447:416], zll_rowround_rowround32_in[415:384], zll_rowround_rowround32_in[383:352], zll_rowround_rowround32_in[127:96], zll_rowround_rowround32_in[351:320], zll_rowround_rowround32_in[319:288], zll_rowround_rowround32_in[287:256], zll_rowround_rowround32_in[255:224], zll_rowround_rowround32_in[223:192], zll_rowround_rowround32_in[191:160], zll_rowround_rowround32_in[159:128], zll_rowround_rowround32_in[95:64], zll_rowround_rowround32_in[63:32], zll_rowround_rowround32_in[31:0]};
  assign zll_rowround_rowround33_in = {zll_rowround_rowround31_in[511:480], zll_rowround_rowround31_in[479:448], zll_rowround_rowround31_in[447:416], zll_rowround_rowround31_in[415:384], zll_rowround_rowround31_in[383:352], zll_rowround_rowround31_in[351:320], zll_rowround_rowround31_in[95:64], zll_rowround_rowround31_in[319:288], zll_rowround_rowround31_in[287:256], zll_rowround_rowround31_in[255:224], zll_rowround_rowround31_in[223:192], zll_rowround_rowround31_in[191:160], zll_rowround_rowround31_in[159:128], zll_rowround_rowround31_in[127:96], zll_rowround_rowround31_in[63:32], zll_rowround_rowround31_in[31:0]};
  assign zll_quarterround_quarterround39_inR5 = {zll_rowround_rowround33_in[255:224], zll_rowround_rowround33_in[479:448], zll_rowround_rowround33_in[511:480], zll_rowround_rowround33_in[415:384]};
  ZLL_QuarterRound_quarterround39  instR5 (zll_quarterround_quarterround39_inR5[127:0], zll_quarterround_quarterround39_outR5);
  assign zll_rowround_rowround25_in = {zll_rowround_rowround33_in[447:416], zll_rowround_rowround33_in[383:352], zll_rowround_rowround33_in[351:320], zll_rowround_rowround33_in[319:288], zll_rowround_rowround33_in[287:256], zll_rowround_rowround33_in[31:0], zll_rowround_rowround33_in[223:192], zll_rowround_rowround33_in[191:160], zll_rowround_rowround33_in[159:128], zll_rowround_rowround33_in[127:96], zll_rowround_rowround33_in[95:64], zll_rowround_rowround33_in[63:32], zll_quarterround_quarterround39_outR5};
  assign zll_rowround_rowround14_in = {zll_rowround_rowround25_in[511:480], zll_rowround_rowround25_in[479:448], zll_rowround_rowround25_in[447:416], zll_rowround_rowround25_in[415:384], zll_rowround_rowround25_in[383:352], zll_rowround_rowround25_in[351:320], zll_rowround_rowround25_in[319:288], zll_rowround_rowround25_in[287:256], zll_rowround_rowround25_in[255:224], zll_rowround_rowround25_in[223:192], zll_rowround_rowround25_in[191:160], zll_rowround_rowround25_in[159:128], zll_rowround_rowround25_in[127:0]};
  assign zll_rowround_rowround7_in = {zll_rowround_rowround14_in[511:480], zll_rowround_rowround14_in[479:448], zll_rowround_rowround14_in[447:416], zll_rowround_rowround14_in[415:384], zll_rowround_rowround14_in[383:352], zll_rowround_rowround14_in[351:320], zll_rowround_rowround14_in[319:288], zll_rowround_rowround14_in[287:256], zll_rowround_rowround14_in[255:224], zll_rowround_rowround14_in[223:192], zll_rowround_rowround14_in[191:160], zll_rowround_rowround14_in[127:96], zll_rowround_rowround14_in[159:128], zll_rowround_rowround14_in[95:64], zll_rowround_rowround14_in[63:32], zll_rowround_rowround14_in[31:0]};
  assign zll_rowround_rowround13_in = {zll_rowround_rowround7_in[511:480], zll_rowround_rowround7_in[95:64], zll_rowround_rowround7_in[479:448], zll_rowround_rowround7_in[447:416], zll_rowround_rowround7_in[415:384], zll_rowround_rowround7_in[383:352], zll_rowround_rowround7_in[351:320], zll_rowround_rowround7_in[319:288], zll_rowround_rowround7_in[287:256], zll_rowround_rowround7_in[255:224], zll_rowround_rowround7_in[223:192], zll_rowround_rowround7_in[191:160], zll_rowround_rowround7_in[159:128], zll_rowround_rowround7_in[127:96], zll_rowround_rowround7_in[63:32], zll_rowround_rowround7_in[31:0]};
  assign zll_rowround_rowround11_in = {zll_rowround_rowround13_in[511:480], zll_rowround_rowround13_in[63:32], zll_rowround_rowround13_in[479:448], zll_rowround_rowround13_in[447:416], zll_rowround_rowround13_in[415:384], zll_rowround_rowround13_in[383:352], zll_rowround_rowround13_in[351:320], zll_rowround_rowround13_in[319:288], zll_rowround_rowround13_in[287:256], zll_rowround_rowround13_in[255:224], zll_rowround_rowround13_in[223:192], zll_rowround_rowround13_in[191:160], zll_rowround_rowround13_in[159:128], zll_rowround_rowround13_in[127:96], zll_rowround_rowround13_in[95:64], zll_rowround_rowround13_in[31:0]};
  assign zll_quarterround_quarterround39_inR6 = {zll_rowround_rowround11_in[223:192], zll_rowround_rowround11_in[191:160], zll_rowround_rowround11_in[159:128], zll_rowround_rowround11_in[511:480]};
  ZLL_QuarterRound_quarterround39  instR6 (zll_quarterround_quarterround39_inR6[127:0], zll_quarterround_quarterround39_outR6);
  assign zll_rowround_rowround2_in = {zll_rowround_rowround11_in[479:448], zll_rowround_rowround11_in[447:416], zll_rowround_rowround11_in[415:384], zll_rowround_rowround11_in[31:0], zll_rowround_rowround11_in[383:352], zll_rowround_rowround11_in[351:320], zll_rowround_rowround11_in[319:288], zll_rowround_rowround11_in[287:256], zll_rowround_rowround11_in[255:224], zll_rowround_rowround11_in[127:96], zll_rowround_rowround11_in[95:64], zll_rowround_rowround11_in[63:32], zll_quarterround_quarterround39_outR6};
  assign zll_rowround_rowround8_in = {zll_rowround_rowround2_in[511:480], zll_rowround_rowround2_in[479:448], zll_rowround_rowround2_in[447:416], zll_rowround_rowround2_in[415:384], zll_rowround_rowround2_in[383:352], zll_rowround_rowround2_in[351:320], zll_rowround_rowround2_in[319:288], zll_rowround_rowround2_in[287:256], zll_rowround_rowround2_in[255:224], zll_rowround_rowround2_in[223:192], zll_rowround_rowround2_in[191:160], zll_rowround_rowround2_in[159:128], zll_rowround_rowround2_in[127:0]};
  assign zll_rowround_rowround12_in = {zll_rowround_rowround8_in[127:96], zll_rowround_rowround8_in[511:480], zll_rowround_rowround8_in[479:448], zll_rowround_rowround8_in[447:416], zll_rowround_rowround8_in[415:384], zll_rowround_rowround8_in[383:352], zll_rowround_rowround8_in[351:320], zll_rowround_rowround8_in[319:288], zll_rowround_rowround8_in[287:256], zll_rowround_rowround8_in[255:224], zll_rowround_rowround8_in[223:192], zll_rowround_rowround8_in[191:160], zll_rowround_rowround8_in[159:128], zll_rowround_rowround8_in[95:64], zll_rowround_rowround8_in[63:32], zll_rowround_rowround8_in[31:0]};
  assign zll_rowround_rowround5_in = {zll_rowround_rowround12_in[511:480], zll_rowround_rowround12_in[479:448], zll_rowround_rowround12_in[447:416], zll_rowround_rowround12_in[415:384], zll_rowround_rowround12_in[383:352], zll_rowround_rowround12_in[351:320], zll_rowround_rowround12_in[319:288], zll_rowround_rowround12_in[287:256], zll_rowround_rowround12_in[255:224], zll_rowround_rowround12_in[95:64], zll_rowround_rowround12_in[223:192], zll_rowround_rowround12_in[191:160], zll_rowround_rowround12_in[159:128], zll_rowround_rowround12_in[127:96], zll_rowround_rowround12_in[63:32], zll_rowround_rowround12_in[31:0]};
  assign zll_rowround_rowround1_in = {zll_rowround_rowround5_in[511:480], zll_rowround_rowround5_in[479:448], zll_rowround_rowround5_in[447:416], zll_rowround_rowround5_in[415:384], zll_rowround_rowround5_in[383:352], zll_rowround_rowround5_in[351:320], zll_rowround_rowround5_in[319:288], zll_rowround_rowround5_in[287:256], zll_rowround_rowround5_in[255:224], zll_rowround_rowround5_in[223:192], zll_rowround_rowround5_in[63:32], zll_rowround_rowround5_in[191:160], zll_rowround_rowround5_in[159:128], zll_rowround_rowround5_in[127:96], zll_rowround_rowround5_in[95:64], zll_rowround_rowround5_in[31:0]};
  assign zll_quarterround_quarterround39_inR7 = {zll_rowround_rowround1_in[415:384], zll_rowround_rowround1_in[159:128], zll_rowround_rowround1_in[127:96], zll_rowround_rowround1_in[287:256]};
  ZLL_QuarterRound_quarterround39  instR7 (zll_quarterround_quarterround39_inR7[127:0], zll_quarterround_quarterround39_outR7);
  assign zll_rowround_rowround21_in = {zll_rowround_rowround1_in[511:480], zll_rowround_rowround1_in[31:0], zll_rowround_rowround1_in[479:448], zll_rowround_rowround1_in[447:416], zll_rowround_rowround1_in[383:352], zll_rowround_rowround1_in[351:320], zll_rowround_rowround1_in[319:288], zll_rowround_rowround1_in[255:224], zll_rowround_rowround1_in[223:192], zll_rowround_rowround1_in[191:160], zll_rowround_rowround1_in[95:64], zll_rowround_rowround1_in[63:32], zll_quarterround_quarterround39_outR7};
  assign zll_rowround_rowround39_in = {zll_rowround_rowround21_in[511:480], zll_rowround_rowround21_in[479:448], zll_rowround_rowround21_in[447:416], zll_rowround_rowround21_in[415:384], zll_rowround_rowround21_in[383:352], zll_rowround_rowround21_in[351:320], zll_rowround_rowround21_in[319:288], zll_rowround_rowround21_in[287:256], zll_rowround_rowround21_in[255:224], zll_rowround_rowround21_in[223:192], zll_rowround_rowround21_in[191:160], zll_rowround_rowround21_in[159:128], zll_rowround_rowround21_in[127:0]};
  assign zll_rowround_rowround27_in = {zll_rowround_rowround39_in[511:480], zll_rowround_rowround39_in[479:448], zll_rowround_rowround39_in[127:96], zll_rowround_rowround39_in[447:416], zll_rowround_rowround39_in[415:384], zll_rowround_rowround39_in[383:352], zll_rowround_rowround39_in[351:320], zll_rowround_rowround39_in[319:288], zll_rowround_rowround39_in[287:256], zll_rowround_rowround39_in[255:224], zll_rowround_rowround39_in[223:192], zll_rowround_rowround39_in[191:160], zll_rowround_rowround39_in[159:128], zll_rowround_rowround39_in[95:64], zll_rowround_rowround39_in[63:32], zll_rowround_rowround39_in[31:0]};
  assign zll_rowround_rowround10_in = {zll_rowround_rowround27_in[95:64], zll_rowround_rowround27_in[511:480], zll_rowround_rowround27_in[479:448], zll_rowround_rowround27_in[447:416], zll_rowround_rowround27_in[415:384], zll_rowround_rowround27_in[383:352], zll_rowround_rowround27_in[351:320], zll_rowround_rowround27_in[319:288], zll_rowround_rowround27_in[287:256], zll_rowround_rowround27_in[255:224], zll_rowround_rowround27_in[223:192], zll_rowround_rowround27_in[191:160], zll_rowround_rowround27_in[159:128], zll_rowround_rowround27_in[127:96], zll_rowround_rowround27_in[63:32], zll_rowround_rowround27_in[31:0]};
  assign lit_in = zll_main_dr12_in[512:0];
  assign res = (lit_in[512] == 1'h0) ? {10'h201{1'h0}} : {1'h1, {zll_rowround_rowround10_in[287:256], zll_rowround_rowround10_in[255:224], zll_rowround_rowround10_in[95:64], zll_rowround_rowround10_in[223:192], zll_rowround_rowround10_in[319:288], zll_rowround_rowround10_in[127:96], zll_rowround_rowround10_in[351:320], zll_rowround_rowround10_in[383:352], zll_rowround_rowround10_in[159:128], zll_rowround_rowround10_in[447:416], zll_rowround_rowround10_in[479:448], zll_rowround_rowround10_in[191:160], zll_rowround_rowround10_in[511:480], zll_rowround_rowround10_in[63:32], zll_rowround_rowround10_in[31:0], zll_rowround_rowround10_in[415:384]}};
endmodule

module Main_conn10 (input logic [5129:0] arg0,
  input logic [512:0] arg1,
  output logic [5129:0] res);
  logic [5642:0] zll_main_conn104_in;
  logic [5642:0] zll_main_conn1010_in;
  logic [5642:0] zll_main_conn1013_in;
  logic [5642:0] zll_main_conn106_in;
  logic [5642:0] zll_main_conn105_in;
  logic [5642:0] zll_main_conn10_in;
  logic [5642:0] zll_main_conn1012_in;
  logic [5129:0] zll_main_conn107_in;
  logic [512:0] main_next_in;
  logic [512:0] main_next_out;
  logic [512:0] main_next_inR1;
  logic [512:0] main_next_outR1;
  logic [512:0] main_next_inR2;
  logic [512:0] main_next_outR2;
  logic [512:0] main_next_inR3;
  logic [512:0] main_next_outR3;
  logic [512:0] main_next_inR4;
  logic [512:0] main_next_outR4;
  logic [512:0] main_next_inR5;
  logic [512:0] main_next_outR5;
  logic [512:0] main_next_inR6;
  logic [512:0] main_next_outR6;
  logic [512:0] main_next_inR7;
  logic [512:0] main_next_outR7;
  logic [512:0] main_next_inR8;
  logic [512:0] main_next_outR8;
  assign zll_main_conn104_in = {arg0, arg1};
  assign zll_main_conn1010_in = zll_main_conn104_in[5642:0];
  assign zll_main_conn1013_in = {zll_main_conn1010_in[5642:5130], zll_main_conn1010_in[4616:4104], zll_main_conn1010_in[5129:4617], zll_main_conn1010_in[4103:3591], zll_main_conn1010_in[3590:3078], zll_main_conn1010_in[3077:2565], zll_main_conn1010_in[2564:2052], zll_main_conn1010_in[2051:1539], zll_main_conn1010_in[1538:1026], zll_main_conn1010_in[1025:513], zll_main_conn1010_in[512:0]};
  assign zll_main_conn106_in = {zll_main_conn1013_in[4103:3591], zll_main_conn1013_in[5642:5130], zll_main_conn1013_in[5129:4617], zll_main_conn1013_in[4616:4104], zll_main_conn1013_in[3590:3078], zll_main_conn1013_in[3077:2565], zll_main_conn1013_in[2564:2052], zll_main_conn1013_in[2051:1539], zll_main_conn1013_in[1538:1026], zll_main_conn1013_in[1025:513], zll_main_conn1013_in[512:0]};
  assign zll_main_conn105_in = {zll_main_conn106_in[5642:5130], zll_main_conn106_in[5129:4617], zll_main_conn106_in[4616:4104], zll_main_conn106_in[3590:3078], zll_main_conn106_in[4103:3591], zll_main_conn106_in[3077:2565], zll_main_conn106_in[2564:2052], zll_main_conn106_in[2051:1539], zll_main_conn106_in[1538:1026], zll_main_conn106_in[1025:513], zll_main_conn106_in[512:0]};
  assign zll_main_conn10_in = {zll_main_conn105_in[2564:2052], zll_main_conn105_in[5642:5130], zll_main_conn105_in[5129:4617], zll_main_conn105_in[4616:4104], zll_main_conn105_in[4103:3591], zll_main_conn105_in[3590:3078], zll_main_conn105_in[3077:2565], zll_main_conn105_in[2051:1539], zll_main_conn105_in[1538:1026], zll_main_conn105_in[1025:513], zll_main_conn105_in[512:0]};
  assign zll_main_conn1012_in = {zll_main_conn10_in[5642:5130], zll_main_conn10_in[5129:4617], zll_main_conn10_in[4616:4104], zll_main_conn10_in[2051:1539], zll_main_conn10_in[4103:3591], zll_main_conn10_in[3590:3078], zll_main_conn10_in[3077:2565], zll_main_conn10_in[2564:2052], zll_main_conn10_in[1538:1026], zll_main_conn10_in[1025:513], zll_main_conn10_in[512:0]};
  assign zll_main_conn107_in = {zll_main_conn1012_in[5642:5130], zll_main_conn1012_in[5129:4617], zll_main_conn1012_in[4616:4104], zll_main_conn1012_in[4103:3591], zll_main_conn1012_in[3590:3078], zll_main_conn1012_in[3077:2565], zll_main_conn1012_in[2564:2052], zll_main_conn1012_in[2051:1539], zll_main_conn1012_in[1538:1026], zll_main_conn1012_in[512:0]};
  assign main_next_in = zll_main_conn107_in[4103:3591];
  Main_next  inst (main_next_in[512:0], main_next_out);
  assign main_next_inR1 = zll_main_conn107_in[2051:1539];
  Main_next  instR1 (main_next_inR1[512:0], main_next_outR1);
  assign main_next_inR2 = zll_main_conn107_in[3077:2565];
  Main_next  instR2 (main_next_inR2[512:0], main_next_outR2);
  assign main_next_inR3 = zll_main_conn107_in[4616:4104];
  Main_next  instR3 (main_next_inR3[512:0], main_next_outR3);
  assign main_next_inR4 = zll_main_conn107_in[2564:2052];
  Main_next  instR4 (main_next_inR4[512:0], main_next_outR4);
  assign main_next_inR5 = zll_main_conn107_in[1538:1026];
  Main_next  instR5 (main_next_inR5[512:0], main_next_outR5);
  assign main_next_inR6 = zll_main_conn107_in[5129:4617];
  Main_next  instR6 (main_next_inR6[512:0], main_next_outR6);
  assign main_next_inR7 = zll_main_conn107_in[3590:3078];
  Main_next  instR7 (main_next_inR7[512:0], main_next_outR7);
  assign main_next_inR8 = zll_main_conn107_in[1025:513];
  Main_next  instR8 (main_next_inR8[512:0], main_next_outR8);
  assign res = {zll_main_conn107_in[512:0], main_next_out, main_next_outR1, main_next_outR2, main_next_outR3, main_next_outR4, main_next_outR5, main_next_outR6, main_next_outR7, main_next_outR8};
endmodule

module Main_next (input logic [512:0] arg0,
  output logic [512:0] res);
  logic [1025:0] zll_main_next1_in;
  logic [512:0] zll_main_next2_in;
  logic [512:0] zll_main_next_in;
  logic [512:0] lit_in;
  assign zll_main_next1_in = {arg0, arg0};
  assign zll_main_next2_in = zll_main_next1_in[1025:513];
  assign zll_main_next_in = zll_main_next2_in[512:0];
  assign lit_in = zll_main_next1_in[512:0];
  assign res = (lit_in[512] == 1'h0) ? {10'h201{1'h0}} : {1'h1, zll_main_next_in[511:0]};
endmodule

module ZLL_Main_out101 (input logic [5129:0] arg0,
  output logic [512:0] res);
  logic [5129:0] zll_main_out102_in;
  logic [4616:0] zll_main_out103_in;
  logic [4103:0] zll_main_out1010_in;
  logic [3590:0] zll_main_out107_in;
  logic [3077:0] zll_main_out105_in;
  logic [2564:0] zll_main_out10_in;
  logic [2051:0] zll_main_out106_in;
  logic [1538:0] zll_main_out104_in;
  logic [1025:0] zll_main_out108_in;
  assign zll_main_out102_in = arg0;
  assign zll_main_out103_in = {zll_main_out102_in[4616:4104], zll_main_out102_in[4103:3591], zll_main_out102_in[3590:3078], zll_main_out102_in[3077:2565], zll_main_out102_in[2564:2052], zll_main_out102_in[2051:1539], zll_main_out102_in[1538:1026], zll_main_out102_in[1025:513], zll_main_out102_in[512:0]};
  assign zll_main_out1010_in = {zll_main_out103_in[4103:3591], zll_main_out103_in[3590:3078], zll_main_out103_in[3077:2565], zll_main_out103_in[2564:2052], zll_main_out103_in[2051:1539], zll_main_out103_in[1538:1026], zll_main_out103_in[1025:513], zll_main_out103_in[512:0]};
  assign zll_main_out107_in = {zll_main_out1010_in[3590:3078], zll_main_out1010_in[3077:2565], zll_main_out1010_in[2564:2052], zll_main_out1010_in[2051:1539], zll_main_out1010_in[1538:1026], zll_main_out1010_in[1025:513], zll_main_out1010_in[512:0]};
  assign zll_main_out105_in = {zll_main_out107_in[3077:2565], zll_main_out107_in[2564:2052], zll_main_out107_in[2051:1539], zll_main_out107_in[1538:1026], zll_main_out107_in[1025:513], zll_main_out107_in[512:0]};
  assign zll_main_out10_in = {zll_main_out105_in[2564:2052], zll_main_out105_in[2051:1539], zll_main_out105_in[1538:1026], zll_main_out105_in[1025:513], zll_main_out105_in[512:0]};
  assign zll_main_out106_in = {zll_main_out10_in[2051:1539], zll_main_out10_in[1538:1026], zll_main_out10_in[1025:513], zll_main_out10_in[512:0]};
  assign zll_main_out104_in = {zll_main_out106_in[1538:1026], zll_main_out106_in[1025:513], zll_main_out106_in[512:0]};
  assign zll_main_out108_in = {zll_main_out104_in[1025:513], zll_main_out104_in[512:0]};
  assign res = zll_main_out108_in[512:0];
endmodule