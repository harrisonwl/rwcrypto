module top_level (input logic [0:0] clk,
  input logic [0:0] rst,
  input logic [0:0] __in0,
  input logic [511:0] __in1,
  output logic [0:0] __out0,
  output logic [511:0] __out1);
  logic [2053:0] zll_pure_dispatch_in;
  logic [1025:0] zll_pure_dispatch4_in;
  logic [1025:0] zll_main_refold1_in;
  logic [1538:0] main_conn21_in;
  logic [1025:0] main_conn21_out;
  logic [1025:0] zll_main_twice3_in;
  logic [1025:0] zll_main_twice3_out;
  logic [1538:0] main_refold1_in;
  logic [2053:0] main_refold1_out;
  logic [2053:0] zll_pure_dispatch5_in;
  logic [512:0] main_refold_in;
  logic [1538:0] main_conn21_inR1;
  logic [1025:0] main_conn21_outR1;
  logic [1025:0] zll_main_twice3_inR1;
  logic [1025:0] zll_main_twice3_outR1;
  logic [1025:0] zll_main_out2_in;
  logic [512:0] zll_main_out2_out;
  logic [2053:0] zll_pure_dispatch2_in;
  logic [2051:0] zll_pure_dispatch1_in;
  logic [2051:0] zll_pure_dispatch3_in;
  logic [2051:0] zll_main_refold_in;
  logic [1538:0] main_conn21_inR2;
  logic [1025:0] main_conn21_outR2;
  logic [1025:0] zll_main_twice3_inR2;
  logic [1025:0] zll_main_twice3_outR2;
  logic [1538:0] main_refold1_inR1;
  logic [2053:0] main_refold1_outR1;
  logic [0:0] __continue;
  logic [1540:0] __resumption_tag;
  logic [1540:0] __resumption_tag_next;
  assign zll_pure_dispatch_in = {{__in0, __in1}, __resumption_tag};
  assign zll_pure_dispatch4_in = {zll_pure_dispatch_in[2053:1541], zll_pure_dispatch_in[512:0]};
  assign zll_main_refold1_in = {zll_pure_dispatch4_in[512:0], zll_pure_dispatch4_in[1025:513]};
  assign main_conn21_in = {{11'h402{1'h0}}, zll_main_refold1_in[1025:513]};
  Main_conn21  inst (main_conn21_in[1538:513], main_conn21_in[512:0], main_conn21_out);
  assign zll_main_twice3_in = main_conn21_out;
  ZLL_Main_twice3  instR1 (zll_main_twice3_in[1025:0], zll_main_twice3_out);
  assign main_refold1_in = {zll_main_twice3_out, zll_main_refold1_in[512:0]};
  Main_refold1  instR2 (main_refold1_in[1538:513], main_refold1_in[512:0], main_refold1_out);
  assign zll_pure_dispatch5_in = {{__in0, __in1}, __resumption_tag};
  assign main_refold_in = zll_pure_dispatch5_in[2053:1541];
  assign main_conn21_inR1 = {{11'h402{1'h0}}, main_refold_in[512:0]};
  Main_conn21  instR3 (main_conn21_inR1[1538:513], main_conn21_inR1[512:0], main_conn21_outR1);
  assign zll_main_twice3_inR1 = main_conn21_outR1;
  ZLL_Main_twice3  instR4 (zll_main_twice3_inR1[1025:0], zll_main_twice3_outR1);
  assign zll_main_out2_in = zll_main_twice3_outR1;
  ZLL_Main_out2  instR5 (zll_main_out2_in[1025:0], zll_main_out2_out);
  assign zll_pure_dispatch2_in = {{__in0, __in1}, __resumption_tag};
  assign zll_pure_dispatch1_in = {zll_pure_dispatch2_in[2053:1541], zll_pure_dispatch2_in[1538:513], zll_pure_dispatch2_in[512:0]};
  assign zll_pure_dispatch3_in = {zll_pure_dispatch1_in[1538:513], zll_pure_dispatch1_in[2051:1539], zll_pure_dispatch1_in[512:0]};
  assign zll_main_refold_in = {zll_pure_dispatch3_in[2051:1026], zll_pure_dispatch3_in[512:0], zll_pure_dispatch3_in[1025:513]};
  assign main_conn21_inR2 = {zll_main_refold_in[2051:1026], zll_main_refold_in[1025:513]};
  Main_conn21  instR6 (main_conn21_inR2[1538:513], main_conn21_inR2[512:0], main_conn21_outR2);
  assign zll_main_twice3_inR2 = main_conn21_outR2;
  ZLL_Main_twice3  instR7 (zll_main_twice3_inR2[1025:0], zll_main_twice3_outR2);
  assign main_refold1_inR1 = {zll_main_twice3_outR2, zll_main_refold_in[512:0]};
  Main_refold1  instR8 (main_refold1_inR1[1538:513], main_refold1_inR1[512:0], main_refold1_outR1);
  assign {__continue, __out0, __out1, __resumption_tag_next} = (zll_pure_dispatch2_in[1540:1539] == 2'h1) ? main_refold1_outR1 : ((zll_pure_dispatch5_in[1540:1539] == 2'h2) ? {zll_main_out2_out, {11'h404{1'h0}}, main_refold_in[512:0]} : main_refold1_out);
  initial __resumption_tag <= {1'h1, {11'h604{1'h0}}};
  always @ (posedge clk or posedge rst) begin
    if (rst == 1'h1) begin
      __resumption_tag <= {1'h1, {11'h604{1'h0}}};
    end else begin
      __resumption_tag <= __resumption_tag_next;
    end
  end
endmodule

module Main_refold1 (input logic [1025:0] arg0,
  input logic [512:0] arg1,
  output logic [2053:0] res);
  logic [1538:0] main_conn21_in;
  logic [1025:0] main_conn21_out;
  logic [1025:0] zll_main_twice3_in;
  logic [1025:0] zll_main_twice3_out;
  logic [1025:0] zll_main_out2_in;
  logic [512:0] zll_main_out2_out;
  assign main_conn21_in = {arg0, arg1};
  Main_conn21  inst (main_conn21_in[1538:513], main_conn21_in[512:0], main_conn21_out);
  assign zll_main_twice3_in = main_conn21_out;
  ZLL_Main_twice3  instR1 (zll_main_twice3_in[1025:0], zll_main_twice3_out);
  assign zll_main_out2_in = zll_main_twice3_out;
  ZLL_Main_out2  instR2 (zll_main_out2_in[1025:0], zll_main_out2_out);
  assign res = {zll_main_out2_out, 2'h1, arg0, arg1};
endmodule

module ZLL_Main_twice3 (input logic [1025:0] arg0,
  output logic [1025:0] res);
  logic [1025:0] zll_main_twice_in;
  logic [512:0] main_io_dr5_in;
  logic [512:0] main_io__dr5_out;
  logic [512:0] main_io_dr5_inR1;
  logic [512:0] main_io__dr5_outR1;
  assign zll_main_twice_in = arg0;
  assign main_io_dr5_in = zll_main_twice_in[1025:513];
  Main_io__dr5  inst (main_io_dr5_in[512:0], main_io__dr5_out);
  assign main_io_dr5_inR1 = zll_main_twice_in[512:0];
  Main_io__dr5  instR1 (main_io_dr5_inR1[512:0], main_io__dr5_outR1);
  assign res = {main_io__dr5_out, main_io__dr5_outR1};
endmodule

module ZLL_ColumnRound_columnround39 (input logic [511:0] arg0,
  output logic [511:0] res);
  logic [511:0] zll_columnround_columnround6_in;
  logic [511:0] zll_columnround_columnround8_in;
  logic [511:0] zll_columnround_columnround34_in;
  logic [511:0] zll_columnround_columnround4_in;
  logic [511:0] zll_columnround_columnround32_in;
  logic [511:0] zll_columnround_columnround12_in;
  logic [511:0] zll_columnround_columnround29_in;
  logic [511:0] zll_columnround_columnround27_in;
  logic [511:0] zll_columnround_columnround36_in;
  logic [511:0] zll_columnround_columnround26_in;
  logic [511:0] zll_columnround_columnround22_in;
  logic [511:0] zll_columnround_columnround5_in;
  logic [511:0] zll_columnround_columnround19_in;
  logic [511:0] zll_columnround_columnround30_in;
  logic [127:0] zll_quarterround_quarterround15_in;
  logic [127:0] zll_quarterround_quarterround15_out;
  logic [511:0] zll_columnround_columnround1_in;
  logic [511:0] zll_columnround_columnround9_in;
  logic [511:0] zll_columnround_columnround11_in;
  logic [511:0] zll_columnround_columnround24_in;
  logic [511:0] zll_columnround_columnround37_in;
  logic [127:0] zll_quarterround_quarterround15_inR1;
  logic [127:0] zll_quarterround_quarterround15_outR1;
  logic [511:0] zll_columnround_columnround7_in;
  logic [511:0] zll_columnround_columnround17_in;
  logic [511:0] zll_columnround_columnround40_in;
  logic [511:0] zll_columnround_columnround25_in;
  logic [511:0] zll_columnround_columnround_in;
  logic [127:0] zll_quarterround_quarterround15_inR2;
  logic [127:0] zll_quarterround_quarterround15_outR2;
  logic [511:0] zll_columnround_columnround16_in;
  logic [511:0] zll_columnround_columnround33_in;
  logic [511:0] zll_columnround_columnround23_in;
  logic [511:0] zll_columnround_columnround31_in;
  logic [511:0] zll_columnround_columnround35_in;
  logic [127:0] zll_quarterround_quarterround15_inR3;
  logic [127:0] zll_quarterround_quarterround15_outR3;
  logic [511:0] zll_columnround_columnround20_in;
  logic [511:0] zll_columnround_columnround38_in;
  logic [511:0] zll_columnround_columnround10_in;
  logic [511:0] zll_columnround_columnround2_in;
  logic [511:0] zll_columnround_columnround18_in;
  assign zll_columnround_columnround6_in = arg0;
  assign zll_columnround_columnround8_in = {zll_columnround_columnround6_in[479:448], zll_columnround_columnround6_in[511:480], zll_columnround_columnround6_in[447:416], zll_columnround_columnround6_in[415:384], zll_columnround_columnround6_in[383:352], zll_columnround_columnround6_in[351:320], zll_columnround_columnround6_in[319:288], zll_columnround_columnround6_in[287:256], zll_columnround_columnround6_in[255:224], zll_columnround_columnround6_in[223:192], zll_columnround_columnround6_in[191:160], zll_columnround_columnround6_in[159:128], zll_columnround_columnround6_in[127:96], zll_columnround_columnround6_in[95:64], zll_columnround_columnround6_in[63:32], zll_columnround_columnround6_in[31:0]};
  assign zll_columnround_columnround34_in = {zll_columnround_columnround8_in[511:480], zll_columnround_columnround8_in[447:416], zll_columnround_columnround8_in[479:448], zll_columnround_columnround8_in[415:384], zll_columnround_columnround8_in[383:352], zll_columnround_columnround8_in[351:320], zll_columnround_columnround8_in[319:288], zll_columnround_columnround8_in[287:256], zll_columnround_columnround8_in[255:224], zll_columnround_columnround8_in[223:192], zll_columnround_columnround8_in[191:160], zll_columnround_columnround8_in[159:128], zll_columnround_columnround8_in[127:96], zll_columnround_columnround8_in[95:64], zll_columnround_columnround8_in[63:32], zll_columnround_columnround8_in[31:0]};
  assign zll_columnround_columnround4_in = {zll_columnround_columnround34_in[511:480], zll_columnround_columnround34_in[479:448], zll_columnround_columnround34_in[415:384], zll_columnround_columnround34_in[447:416], zll_columnround_columnround34_in[383:352], zll_columnround_columnround34_in[351:320], zll_columnround_columnround34_in[319:288], zll_columnround_columnround34_in[287:256], zll_columnround_columnround34_in[255:224], zll_columnround_columnround34_in[223:192], zll_columnround_columnround34_in[191:160], zll_columnround_columnround34_in[159:128], zll_columnround_columnround34_in[127:96], zll_columnround_columnround34_in[95:64], zll_columnround_columnround34_in[63:32], zll_columnround_columnround34_in[31:0]};
  assign zll_columnround_columnround32_in = {zll_columnround_columnround4_in[351:320], zll_columnround_columnround4_in[511:480], zll_columnround_columnround4_in[479:448], zll_columnround_columnround4_in[447:416], zll_columnround_columnround4_in[415:384], zll_columnround_columnround4_in[383:352], zll_columnround_columnround4_in[319:288], zll_columnround_columnround4_in[287:256], zll_columnround_columnround4_in[255:224], zll_columnround_columnround4_in[223:192], zll_columnround_columnround4_in[191:160], zll_columnround_columnround4_in[159:128], zll_columnround_columnround4_in[127:96], zll_columnround_columnround4_in[95:64], zll_columnround_columnround4_in[63:32], zll_columnround_columnround4_in[31:0]};
  assign zll_columnround_columnround12_in = {zll_columnround_columnround32_in[511:480], zll_columnround_columnround32_in[479:448], zll_columnround_columnround32_in[319:288], zll_columnround_columnround32_in[447:416], zll_columnround_columnround32_in[415:384], zll_columnround_columnround32_in[383:352], zll_columnround_columnround32_in[351:320], zll_columnround_columnround32_in[287:256], zll_columnround_columnround32_in[255:224], zll_columnround_columnround32_in[223:192], zll_columnround_columnround32_in[191:160], zll_columnround_columnround32_in[159:128], zll_columnround_columnround32_in[127:96], zll_columnround_columnround32_in[95:64], zll_columnround_columnround32_in[63:32], zll_columnround_columnround32_in[31:0]};
  assign zll_columnround_columnround29_in = {zll_columnround_columnround12_in[511:480], zll_columnround_columnround12_in[479:448], zll_columnround_columnround12_in[447:416], zll_columnround_columnround12_in[415:384], zll_columnround_columnround12_in[383:352], zll_columnround_columnround12_in[287:256], zll_columnround_columnround12_in[351:320], zll_columnround_columnround12_in[319:288], zll_columnround_columnround12_in[255:224], zll_columnround_columnround12_in[223:192], zll_columnround_columnround12_in[191:160], zll_columnround_columnround12_in[159:128], zll_columnround_columnround12_in[127:96], zll_columnround_columnround12_in[95:64], zll_columnround_columnround12_in[63:32], zll_columnround_columnround12_in[31:0]};
  assign zll_columnround_columnround27_in = {zll_columnround_columnround29_in[511:480], zll_columnround_columnround29_in[479:448], zll_columnround_columnround29_in[447:416], zll_columnround_columnround29_in[415:384], zll_columnround_columnround29_in[383:352], zll_columnround_columnround29_in[255:224], zll_columnround_columnround29_in[351:320], zll_columnround_columnround29_in[319:288], zll_columnround_columnround29_in[287:256], zll_columnround_columnround29_in[223:192], zll_columnround_columnround29_in[191:160], zll_columnround_columnround29_in[159:128], zll_columnround_columnround29_in[127:96], zll_columnround_columnround29_in[95:64], zll_columnround_columnround29_in[63:32], zll_columnround_columnround29_in[31:0]};
  assign zll_columnround_columnround36_in = {zll_columnround_columnround27_in[511:480], zll_columnround_columnround27_in[479:448], zll_columnround_columnround27_in[447:416], zll_columnround_columnround27_in[415:384], zll_columnround_columnround27_in[383:352], zll_columnround_columnround27_in[351:320], zll_columnround_columnround27_in[319:288], zll_columnround_columnround27_in[223:192], zll_columnround_columnround27_in[287:256], zll_columnround_columnround27_in[255:224], zll_columnround_columnround27_in[191:160], zll_columnround_columnround27_in[159:128], zll_columnround_columnround27_in[127:96], zll_columnround_columnround27_in[95:64], zll_columnround_columnround27_in[63:32], zll_columnround_columnround27_in[31:0]};
  assign zll_columnround_columnround26_in = {zll_columnround_columnround36_in[511:480], zll_columnround_columnround36_in[479:448], zll_columnround_columnround36_in[447:416], zll_columnround_columnround36_in[191:160], zll_columnround_columnround36_in[415:384], zll_columnround_columnround36_in[383:352], zll_columnround_columnround36_in[351:320], zll_columnround_columnround36_in[319:288], zll_columnround_columnround36_in[287:256], zll_columnround_columnround36_in[255:224], zll_columnround_columnround36_in[223:192], zll_columnround_columnround36_in[159:128], zll_columnround_columnround36_in[127:96], zll_columnround_columnround36_in[95:64], zll_columnround_columnround36_in[63:32], zll_columnround_columnround36_in[31:0]};
  assign zll_columnround_columnround22_in = {zll_columnround_columnround26_in[511:480], zll_columnround_columnround26_in[479:448], zll_columnround_columnround26_in[447:416], zll_columnround_columnround26_in[415:384], zll_columnround_columnround26_in[383:352], zll_columnround_columnround26_in[159:128], zll_columnround_columnround26_in[351:320], zll_columnround_columnround26_in[319:288], zll_columnround_columnround26_in[287:256], zll_columnround_columnround26_in[255:224], zll_columnround_columnround26_in[223:192], zll_columnround_columnround26_in[191:160], zll_columnround_columnround26_in[127:96], zll_columnround_columnround26_in[95:64], zll_columnround_columnround26_in[63:32], zll_columnround_columnround26_in[31:0]};
  assign zll_columnround_columnround5_in = {zll_columnround_columnround22_in[127:96], zll_columnround_columnround22_in[511:480], zll_columnround_columnround22_in[479:448], zll_columnround_columnround22_in[447:416], zll_columnround_columnround22_in[415:384], zll_columnround_columnround22_in[383:352], zll_columnround_columnround22_in[351:320], zll_columnround_columnround22_in[319:288], zll_columnround_columnround22_in[287:256], zll_columnround_columnround22_in[255:224], zll_columnround_columnround22_in[223:192], zll_columnround_columnround22_in[191:160], zll_columnround_columnround22_in[159:128], zll_columnround_columnround22_in[95:64], zll_columnround_columnround22_in[63:32], zll_columnround_columnround22_in[31:0]};
  assign zll_columnround_columnround19_in = {zll_columnround_columnround5_in[511:480], zll_columnround_columnround5_in[479:448], zll_columnround_columnround5_in[447:416], zll_columnround_columnround5_in[415:384], zll_columnround_columnround5_in[383:352], zll_columnround_columnround5_in[351:320], zll_columnround_columnround5_in[319:288], zll_columnround_columnround5_in[287:256], zll_columnround_columnround5_in[95:64], zll_columnround_columnround5_in[255:224], zll_columnround_columnround5_in[223:192], zll_columnround_columnround5_in[191:160], zll_columnround_columnround5_in[159:128], zll_columnround_columnround5_in[127:96], zll_columnround_columnround5_in[63:32], zll_columnround_columnround5_in[31:0]};
  assign zll_columnround_columnround30_in = {zll_columnround_columnround19_in[511:480], zll_columnround_columnround19_in[479:448], zll_columnround_columnround19_in[447:416], zll_columnround_columnround19_in[415:384], zll_columnround_columnround19_in[383:352], zll_columnround_columnround19_in[351:320], zll_columnround_columnround19_in[319:288], zll_columnround_columnround19_in[287:256], zll_columnround_columnround19_in[255:224], zll_columnround_columnround19_in[223:192], zll_columnround_columnround19_in[63:32], zll_columnround_columnround19_in[191:160], zll_columnround_columnround19_in[159:128], zll_columnround_columnround19_in[127:96], zll_columnround_columnround19_in[95:64], zll_columnround_columnround19_in[31:0]};
  assign zll_quarterround_quarterround15_in = {zll_columnround_columnround30_in[95:64], zll_columnround_columnround30_in[63:32], zll_columnround_columnround30_in[223:192], zll_columnround_columnround30_in[511:480]};
  ZLL_QuarterRound_quarterround15  inst (zll_quarterround_quarterround15_in[127:0], zll_quarterround_quarterround15_out);
  assign zll_columnround_columnround1_in = {zll_columnround_columnround30_in[479:448], zll_columnround_columnround30_in[447:416], zll_columnround_columnround30_in[415:384], zll_columnround_columnround30_in[31:0], zll_columnround_columnround30_in[383:352], zll_columnround_columnround30_in[351:320], zll_columnround_columnround30_in[319:288], zll_columnround_columnround30_in[287:256], zll_columnround_columnround30_in[255:224], zll_columnround_columnround30_in[191:160], zll_columnround_columnround30_in[159:128], zll_columnround_columnround30_in[127:96], zll_quarterround_quarterround15_out};
  assign zll_columnround_columnround9_in = {zll_columnround_columnround1_in[511:480], zll_columnround_columnround1_in[479:448], zll_columnround_columnround1_in[447:416], zll_columnround_columnround1_in[415:384], zll_columnround_columnround1_in[383:352], zll_columnround_columnround1_in[351:320], zll_columnround_columnround1_in[319:288], zll_columnround_columnround1_in[287:256], zll_columnround_columnround1_in[255:224], zll_columnround_columnround1_in[223:192], zll_columnround_columnround1_in[191:160], zll_columnround_columnround1_in[159:128], zll_columnround_columnround1_in[127:0]};
  assign zll_columnround_columnround11_in = {zll_columnround_columnround9_in[511:480], zll_columnround_columnround9_in[479:448], zll_columnround_columnround9_in[447:416], zll_columnround_columnround9_in[415:384], zll_columnround_columnround9_in[383:352], zll_columnround_columnround9_in[351:320], zll_columnround_columnround9_in[319:288], zll_columnround_columnround9_in[287:256], zll_columnround_columnround9_in[255:224], zll_columnround_columnround9_in[223:192], zll_columnround_columnround9_in[127:96], zll_columnround_columnround9_in[191:160], zll_columnround_columnround9_in[159:128], zll_columnround_columnround9_in[95:64], zll_columnround_columnround9_in[63:32], zll_columnround_columnround9_in[31:0]};
  assign zll_columnround_columnround24_in = {zll_columnround_columnround11_in[511:480], zll_columnround_columnround11_in[479:448], zll_columnround_columnround11_in[447:416], zll_columnround_columnround11_in[415:384], zll_columnround_columnround11_in[383:352], zll_columnround_columnround11_in[351:320], zll_columnround_columnround11_in[319:288], zll_columnround_columnround11_in[287:256], zll_columnround_columnround11_in[255:224], zll_columnround_columnround11_in[223:192], zll_columnround_columnround11_in[95:64], zll_columnround_columnround11_in[191:160], zll_columnround_columnround11_in[159:128], zll_columnround_columnround11_in[127:96], zll_columnround_columnround11_in[63:32], zll_columnround_columnround11_in[31:0]};
  assign zll_columnround_columnround37_in = {zll_columnround_columnround24_in[511:480], zll_columnround_columnround24_in[479:448], zll_columnround_columnround24_in[447:416], zll_columnround_columnround24_in[415:384], zll_columnround_columnround24_in[383:352], zll_columnround_columnround24_in[351:320], zll_columnround_columnround24_in[319:288], zll_columnround_columnround24_in[63:32], zll_columnround_columnround24_in[287:256], zll_columnround_columnround24_in[255:224], zll_columnround_columnround24_in[223:192], zll_columnround_columnround24_in[191:160], zll_columnround_columnround24_in[159:128], zll_columnround_columnround24_in[127:96], zll_columnround_columnround24_in[95:64], zll_columnround_columnround24_in[31:0]};
  assign zll_quarterround_quarterround15_inR1 = {zll_columnround_columnround37_in[511:480], zll_columnround_columnround37_in[63:32], zll_columnround_columnround37_in[223:192], zll_columnround_columnround37_in[479:448]};
  ZLL_QuarterRound_quarterround15  instR1 (zll_quarterround_quarterround15_inR1[127:0], zll_quarterround_quarterround15_outR1);
  assign zll_columnround_columnround7_in = {zll_columnround_columnround37_in[31:0], zll_columnround_columnround37_in[447:416], zll_columnround_columnround37_in[415:384], zll_columnround_columnround37_in[383:352], zll_columnround_columnround37_in[351:320], zll_columnround_columnround37_in[319:288], zll_columnround_columnround37_in[287:256], zll_columnround_columnround37_in[255:224], zll_columnround_columnround37_in[191:160], zll_columnround_columnround37_in[159:128], zll_columnround_columnround37_in[127:96], zll_columnround_columnround37_in[95:64], zll_quarterround_quarterround15_outR1};
  assign zll_columnround_columnround17_in = {zll_columnround_columnround7_in[511:480], zll_columnround_columnround7_in[479:448], zll_columnround_columnround7_in[447:416], zll_columnround_columnround7_in[415:384], zll_columnround_columnround7_in[383:352], zll_columnround_columnround7_in[351:320], zll_columnround_columnround7_in[319:288], zll_columnround_columnround7_in[287:256], zll_columnround_columnround7_in[255:224], zll_columnround_columnround7_in[223:192], zll_columnround_columnround7_in[191:160], zll_columnround_columnround7_in[159:128], zll_columnround_columnround7_in[127:0]};
  assign zll_columnround_columnround40_in = {zll_columnround_columnround17_in[127:96], zll_columnround_columnround17_in[511:480], zll_columnround_columnround17_in[479:448], zll_columnround_columnround17_in[447:416], zll_columnround_columnround17_in[415:384], zll_columnround_columnround17_in[383:352], zll_columnround_columnround17_in[351:320], zll_columnround_columnround17_in[319:288], zll_columnround_columnround17_in[287:256], zll_columnround_columnround17_in[255:224], zll_columnround_columnround17_in[223:192], zll_columnround_columnround17_in[191:160], zll_columnround_columnround17_in[159:128], zll_columnround_columnround17_in[95:64], zll_columnround_columnround17_in[63:32], zll_columnround_columnround17_in[31:0]};
  assign zll_columnround_columnround25_in = {zll_columnround_columnround40_in[511:480], zll_columnround_columnround40_in[479:448], zll_columnround_columnround40_in[447:416], zll_columnround_columnround40_in[415:384], zll_columnround_columnround40_in[383:352], zll_columnround_columnround40_in[351:320], zll_columnround_columnround40_in[319:288], zll_columnround_columnround40_in[287:256], zll_columnround_columnround40_in[255:224], zll_columnround_columnround40_in[223:192], zll_columnround_columnround40_in[95:64], zll_columnround_columnround40_in[191:160], zll_columnround_columnround40_in[159:128], zll_columnround_columnround40_in[127:96], zll_columnround_columnround40_in[63:32], zll_columnround_columnround40_in[31:0]};
  assign zll_columnround_columnround_in = {zll_columnround_columnround25_in[511:480], zll_columnround_columnround25_in[479:448], zll_columnround_columnround25_in[447:416], zll_columnround_columnround25_in[415:384], zll_columnround_columnround25_in[383:352], zll_columnround_columnround25_in[351:320], zll_columnround_columnround25_in[319:288], zll_columnround_columnround25_in[287:256], zll_columnround_columnround25_in[255:224], zll_columnround_columnround25_in[63:32], zll_columnround_columnround25_in[223:192], zll_columnround_columnround25_in[191:160], zll_columnround_columnround25_in[159:128], zll_columnround_columnround25_in[127:96], zll_columnround_columnround25_in[95:64], zll_columnround_columnround25_in[31:0]};
  assign zll_quarterround_quarterround15_inR2 = {zll_columnround_columnround_in[383:352], zll_columnround_columnround_in[191:160], zll_columnround_columnround_in[351:320], zll_columnround_columnround_in[447:416]};
  ZLL_QuarterRound_quarterround15  instR2 (zll_quarterround_quarterround15_inR2[127:0], zll_quarterround_quarterround15_outR2);
  assign zll_columnround_columnround16_in = {zll_columnround_columnround_in[31:0], zll_columnround_columnround_in[511:480], zll_columnround_columnround_in[479:448], zll_columnround_columnround_in[415:384], zll_columnround_columnround_in[319:288], zll_columnround_columnround_in[287:256], zll_columnround_columnround_in[255:224], zll_columnround_columnround_in[223:192], zll_columnround_columnround_in[159:128], zll_columnround_columnround_in[127:96], zll_columnround_columnround_in[95:64], zll_columnround_columnround_in[63:32], zll_quarterround_quarterround15_outR2};
  assign zll_columnround_columnround33_in = {zll_columnround_columnround16_in[511:480], zll_columnround_columnround16_in[479:448], zll_columnround_columnround16_in[447:416], zll_columnround_columnround16_in[415:384], zll_columnround_columnround16_in[383:352], zll_columnround_columnround16_in[351:320], zll_columnround_columnround16_in[319:288], zll_columnround_columnround16_in[287:256], zll_columnround_columnround16_in[255:224], zll_columnround_columnround16_in[223:192], zll_columnround_columnround16_in[191:160], zll_columnround_columnround16_in[159:128], zll_columnround_columnround16_in[127:0]};
  assign zll_columnround_columnround23_in = {zll_columnround_columnround33_in[511:480], zll_columnround_columnround33_in[479:448], zll_columnround_columnround33_in[447:416], zll_columnround_columnround33_in[415:384], zll_columnround_columnround33_in[127:96], zll_columnround_columnround33_in[383:352], zll_columnround_columnround33_in[351:320], zll_columnround_columnround33_in[319:288], zll_columnround_columnround33_in[287:256], zll_columnround_columnround33_in[255:224], zll_columnround_columnround33_in[223:192], zll_columnround_columnround33_in[191:160], zll_columnround_columnround33_in[159:128], zll_columnround_columnround33_in[95:64], zll_columnround_columnround33_in[63:32], zll_columnround_columnround33_in[31:0]};
  assign zll_columnround_columnround31_in = {zll_columnround_columnround23_in[511:480], zll_columnround_columnround23_in[479:448], zll_columnround_columnround23_in[95:64], zll_columnround_columnround23_in[447:416], zll_columnround_columnround23_in[415:384], zll_columnround_columnround23_in[383:352], zll_columnround_columnround23_in[351:320], zll_columnround_columnround23_in[319:288], zll_columnround_columnround23_in[287:256], zll_columnround_columnround23_in[255:224], zll_columnround_columnround23_in[223:192], zll_columnround_columnround23_in[191:160], zll_columnround_columnround23_in[159:128], zll_columnround_columnround23_in[127:96], zll_columnround_columnround23_in[63:32], zll_columnround_columnround23_in[31:0]};
  assign zll_columnround_columnround35_in = {zll_columnround_columnround31_in[511:480], zll_columnround_columnround31_in[479:448], zll_columnround_columnround31_in[447:416], zll_columnround_columnround31_in[415:384], zll_columnround_columnround31_in[383:352], zll_columnround_columnround31_in[351:320], zll_columnround_columnround31_in[319:288], zll_columnround_columnround31_in[287:256], zll_columnround_columnround31_in[255:224], zll_columnround_columnround31_in[63:32], zll_columnround_columnround31_in[223:192], zll_columnround_columnround31_in[191:160], zll_columnround_columnround31_in[159:128], zll_columnround_columnround31_in[127:96], zll_columnround_columnround31_in[95:64], zll_columnround_columnround31_in[31:0]};
  assign zll_quarterround_quarterround15_inR3 = {zll_columnround_columnround35_in[383:352], zll_columnround_columnround35_in[255:224], zll_columnround_columnround35_in[63:32], zll_columnround_columnround35_in[319:288]};
  ZLL_QuarterRound_quarterround15  instR3 (zll_quarterround_quarterround15_inR3[127:0], zll_quarterround_quarterround15_outR3);
  assign zll_columnround_columnround20_in = {zll_columnround_columnround35_in[511:480], zll_columnround_columnround35_in[479:448], zll_columnround_columnround35_in[447:416], zll_columnround_columnround35_in[415:384], zll_columnround_columnround35_in[351:320], zll_columnround_columnround35_in[287:256], zll_columnround_columnround35_in[223:192], zll_columnround_columnround35_in[191:160], zll_columnround_columnround35_in[159:128], zll_columnround_columnround35_in[127:96], zll_columnround_columnround35_in[31:0], zll_columnround_columnround35_in[95:64], zll_quarterround_quarterround15_outR3};
  assign zll_columnround_columnround38_in = {zll_columnround_columnround20_in[511:480], zll_columnround_columnround20_in[479:448], zll_columnround_columnround20_in[447:416], zll_columnround_columnround20_in[415:384], zll_columnround_columnround20_in[383:352], zll_columnround_columnround20_in[351:320], zll_columnround_columnround20_in[319:288], zll_columnround_columnround20_in[287:256], zll_columnround_columnround20_in[255:224], zll_columnround_columnround20_in[223:192], zll_columnround_columnround20_in[191:160], zll_columnround_columnround20_in[159:128], zll_columnround_columnround20_in[127:0]};
  assign zll_columnround_columnround10_in = {zll_columnround_columnround38_in[511:480], zll_columnround_columnround38_in[479:448], zll_columnround_columnround38_in[447:416], zll_columnround_columnround38_in[415:384], zll_columnround_columnround38_in[127:96], zll_columnround_columnround38_in[383:352], zll_columnround_columnround38_in[351:320], zll_columnround_columnround38_in[319:288], zll_columnround_columnround38_in[287:256], zll_columnround_columnround38_in[255:224], zll_columnround_columnround38_in[223:192], zll_columnround_columnround38_in[191:160], zll_columnround_columnround38_in[159:128], zll_columnround_columnround38_in[95:64], zll_columnround_columnround38_in[63:32], zll_columnround_columnround38_in[31:0]};
  assign zll_columnround_columnround2_in = {zll_columnround_columnround10_in[511:480], zll_columnround_columnround10_in[479:448], zll_columnround_columnround10_in[447:416], zll_columnround_columnround10_in[415:384], zll_columnround_columnround10_in[383:352], zll_columnround_columnround10_in[95:64], zll_columnround_columnround10_in[351:320], zll_columnround_columnround10_in[319:288], zll_columnround_columnround10_in[287:256], zll_columnround_columnround10_in[255:224], zll_columnround_columnround10_in[223:192], zll_columnround_columnround10_in[191:160], zll_columnround_columnround10_in[159:128], zll_columnround_columnround10_in[127:96], zll_columnround_columnround10_in[63:32], zll_columnround_columnround10_in[31:0]};
  assign zll_columnround_columnround18_in = {zll_columnround_columnround2_in[63:32], zll_columnround_columnround2_in[511:480], zll_columnround_columnround2_in[479:448], zll_columnround_columnround2_in[447:416], zll_columnround_columnround2_in[415:384], zll_columnround_columnround2_in[383:352], zll_columnround_columnround2_in[351:320], zll_columnround_columnround2_in[319:288], zll_columnround_columnround2_in[287:256], zll_columnround_columnround2_in[255:224], zll_columnround_columnround2_in[223:192], zll_columnround_columnround2_in[191:160], zll_columnround_columnround2_in[159:128], zll_columnround_columnround2_in[127:96], zll_columnround_columnround2_in[95:64], zll_columnround_columnround2_in[31:0]};
  assign res = {zll_columnround_columnround18_in[63:32], zll_columnround_columnround18_in[479:448], zll_columnround_columnround18_in[223:192], zll_columnround_columnround18_in[319:288], zll_columnround_columnround18_in[127:96], zll_columnround_columnround18_in[447:416], zll_columnround_columnround18_in[95:64], zll_columnround_columnround18_in[511:480], zll_columnround_columnround18_in[255:224], zll_columnround_columnround18_in[159:128], zll_columnround_columnround18_in[287:256], zll_columnround_columnround18_in[31:0], zll_columnround_columnround18_in[383:352], zll_columnround_columnround18_in[191:160], zll_columnround_columnround18_in[415:384], zll_columnround_columnround18_in[351:320]};
endmodule

module Main_conn21 (input logic [1025:0] arg0,
  input logic [512:0] arg1,
  output logic [1025:0] res);
  logic [1538:0] zll_main_conn24_in;
  logic [1538:0] zll_main_conn2_in;
  logic [1025:0] zll_main_conn21_in;
  logic [512:0] main_next_in;
  logic [1025:0] zll_main_next1_in;
  logic [512:0] zll_main_next_in;
  logic [512:0] zll_main_next2_in;
  logic [512:0] lit_in;
  assign zll_main_conn24_in = {arg0, arg1};
  assign zll_main_conn2_in = zll_main_conn24_in[1538:0];
  assign zll_main_conn21_in = {zll_main_conn2_in[1538:1026], zll_main_conn2_in[512:0]};
  assign main_next_in = zll_main_conn21_in[1025:513];
  assign zll_main_next1_in = {main_next_in[512:0], main_next_in[512:0]};
  assign zll_main_next_in = zll_main_next1_in[1025:513];
  assign zll_main_next2_in = zll_main_next_in[512:0];
  assign lit_in = zll_main_next1_in[512:0];
  assign res = {zll_main_conn21_in[512:0], (lit_in[512] == 1'h0) ? {10'h201{1'h0}} : {1'h1, zll_main_next2_in[511:0]}};
endmodule

module ZLL_QuarterRound_quarterround32 (input logic [63:0] arg0,
  output logic [31:0] res);
  logic [63:0] zll_quarterround_quarterround20_in;
  logic [63:0] binop_in;
  logic [63:0] binop_inR1;
  logic [63:0] binop_inR2;
  logic [63:0] binop_inR3;
  assign zll_quarterround_quarterround20_in = arg0;
  assign binop_in = {zll_quarterround_quarterround20_in[31:0], zll_quarterround_quarterround20_in[63:32]};
  assign binop_inR1 = {32'h20, zll_quarterround_quarterround20_in[63:32]};
  assign binop_inR2 = {zll_quarterround_quarterround20_in[31:0], binop_inR1[63:32] - binop_inR1[31:0]};
  assign binop_inR3 = {binop_in[63:32] << binop_in[31:0], binop_inR2[63:32] >> binop_inR2[31:0]};
  assign res = binop_inR3[63:32] | binop_inR3[31:0];
endmodule

module ZLL_QuarterRound_quarterround15 (input logic [127:0] arg0,
  output logic [127:0] res);
  logic [127:0] zll_quarterround_quarterround38_in;
  logic [63:0] binop_in;
  logic [31:0] zll_quarterround_quarterround35_in;
  logic [63:0] zll_quarterround_quarterround32_in;
  logic [31:0] zll_quarterround_quarterround32_out;
  logic [63:0] binop_inR1;
  logic [127:0] zll_quarterround_quarterround_in;
  logic [63:0] binop_inR2;
  logic [31:0] zll_quarterround_quarterround8_in;
  logic [63:0] zll_quarterround_quarterround32_inR1;
  logic [31:0] zll_quarterround_quarterround32_outR1;
  logic [63:0] binop_inR3;
  logic [127:0] zll_quarterround_quarterround26_in;
  logic [63:0] binop_inR4;
  logic [31:0] zll_quarterround_quarterround17_in;
  logic [63:0] zll_quarterround_quarterround32_inR2;
  logic [31:0] zll_quarterround_quarterround32_outR2;
  logic [63:0] binop_inR5;
  logic [127:0] zll_quarterround_quarterround19_in;
  logic [63:0] binop_inR6;
  logic [31:0] zll_quarterround_quarterround37_in;
  logic [63:0] zll_quarterround_quarterround32_inR3;
  logic [31:0] zll_quarterround_quarterround32_outR3;
  logic [63:0] binop_inR7;
  logic [127:0] zll_quarterround_quarterround3_in;
  assign zll_quarterround_quarterround38_in = arg0;
  assign binop_in = {zll_quarterround_quarterround38_in[127:96], zll_quarterround_quarterround38_in[31:0]};
  assign zll_quarterround_quarterround35_in = binop_in[63:32] + binop_in[31:0];
  assign zll_quarterround_quarterround32_in = {32'h7, zll_quarterround_quarterround35_in[31:0]};
  ZLL_QuarterRound_quarterround32  inst (zll_quarterround_quarterround32_in[63:0], zll_quarterround_quarterround32_out);
  assign binop_inR1 = {zll_quarterround_quarterround38_in[95:64], zll_quarterround_quarterround32_out};
  assign zll_quarterround_quarterround_in = {zll_quarterround_quarterround38_in[127:96], zll_quarterround_quarterround38_in[63:32], zll_quarterround_quarterround38_in[31:0], binop_inR1[63:32] ^ binop_inR1[31:0]};
  assign binop_inR2 = {zll_quarterround_quarterround_in[31:0], zll_quarterround_quarterround_in[127:96]};
  assign zll_quarterround_quarterround8_in = binop_inR2[63:32] + binop_inR2[31:0];
  assign zll_quarterround_quarterround32_inR1 = {32'h9, zll_quarterround_quarterround8_in[31:0]};
  ZLL_QuarterRound_quarterround32  instR1 (zll_quarterround_quarterround32_inR1[63:0], zll_quarterround_quarterround32_outR1);
  assign binop_inR3 = {zll_quarterround_quarterround_in[95:64], zll_quarterround_quarterround32_outR1};
  assign zll_quarterround_quarterround26_in = {zll_quarterround_quarterround_in[127:96], zll_quarterround_quarterround_in[31:0], zll_quarterround_quarterround_in[63:32], binop_inR3[63:32] ^ binop_inR3[31:0]};
  assign binop_inR4 = {zll_quarterround_quarterround26_in[31:0], zll_quarterround_quarterround26_in[95:64]};
  assign zll_quarterround_quarterround17_in = binop_inR4[63:32] + binop_inR4[31:0];
  assign zll_quarterround_quarterround32_inR2 = {32'hd, zll_quarterround_quarterround17_in[31:0]};
  ZLL_QuarterRound_quarterround32  instR2 (zll_quarterround_quarterround32_inR2[63:0], zll_quarterround_quarterround32_outR2);
  assign binop_inR5 = {zll_quarterround_quarterround26_in[63:32], zll_quarterround_quarterround32_outR2};
  assign zll_quarterround_quarterround19_in = {zll_quarterround_quarterround26_in[127:96], zll_quarterround_quarterround26_in[31:0], zll_quarterround_quarterround26_in[95:64], binop_inR5[63:32] ^ binop_inR5[31:0]};
  assign binop_inR6 = {zll_quarterround_quarterround19_in[31:0], zll_quarterround_quarterround19_in[95:64]};
  assign zll_quarterround_quarterround37_in = binop_inR6[63:32] + binop_inR6[31:0];
  assign zll_quarterround_quarterround32_inR3 = {32'h12, zll_quarterround_quarterround37_in[31:0]};
  ZLL_QuarterRound_quarterround32  instR3 (zll_quarterround_quarterround32_inR3[63:0], zll_quarterround_quarterround32_outR3);
  assign binop_inR7 = {zll_quarterround_quarterround19_in[127:96], zll_quarterround_quarterround32_outR3};
  assign zll_quarterround_quarterround3_in = {zll_quarterround_quarterround19_in[95:64], zll_quarterround_quarterround19_in[63:32], zll_quarterround_quarterround19_in[31:0], binop_inR7[63:32] ^ binop_inR7[31:0]};
  assign res = {zll_quarterround_quarterround3_in[31:0], zll_quarterround_quarterround3_in[95:64], zll_quarterround_quarterround3_in[127:96], zll_quarterround_quarterround3_in[63:32]};
endmodule

module Main_io__dr5 (input logic [512:0] arg0,
  output logic [512:0] res);
  logic [1025:0] zll_main_io_dr51_in;
  logic [512:0] zll_main_io_dr5_in;
  logic [512:0] zll_main_io_dr53_in;
  logic [511:0] zll_columnround_columnround39_in;
  logic [511:0] zll_columnround_columnround39_out;
  logic [511:0] zll_rowround_rowround10_in;
  logic [511:0] zll_rowround_rowround10_out;
  logic [511:0] zll_columnround_columnround39_inR1;
  logic [511:0] zll_columnround_columnround39_outR1;
  logic [511:0] zll_rowround_rowround10_inR1;
  logic [511:0] zll_rowround_rowround10_outR1;
  logic [511:0] zll_columnround_columnround39_inR2;
  logic [511:0] zll_columnround_columnround39_outR2;
  logic [511:0] zll_rowround_rowround10_inR2;
  logic [511:0] zll_rowround_rowround10_outR2;
  logic [511:0] zll_columnround_columnround39_inR3;
  logic [511:0] zll_columnround_columnround39_outR3;
  logic [511:0] zll_rowround_rowround10_inR3;
  logic [511:0] zll_rowround_rowround10_outR3;
  logic [511:0] zll_columnround_columnround39_inR4;
  logic [511:0] zll_columnround_columnround39_outR4;
  logic [511:0] zll_rowround_rowround10_inR4;
  logic [511:0] zll_rowround_rowround10_outR4;
  logic [512:0] lit_in;
  assign zll_main_io_dr51_in = {arg0, arg0};
  assign zll_main_io_dr5_in = zll_main_io_dr51_in[1025:513];
  assign zll_main_io_dr53_in = zll_main_io_dr5_in[512:0];
  assign zll_columnround_columnround39_in = zll_main_io_dr53_in[511:0];
  ZLL_ColumnRound_columnround39  inst (zll_columnround_columnround39_in[511:0], zll_columnround_columnround39_out);
  assign zll_rowround_rowround10_in = zll_columnround_columnround39_out;
  ZLL_RowRound_rowround10  instR1 (zll_rowround_rowround10_in[511:0], zll_rowround_rowround10_out);
  assign zll_columnround_columnround39_inR1 = zll_rowround_rowround10_out;
  ZLL_ColumnRound_columnround39  instR2 (zll_columnround_columnround39_inR1[511:0], zll_columnround_columnround39_outR1);
  assign zll_rowround_rowround10_inR1 = zll_columnround_columnround39_outR1;
  ZLL_RowRound_rowround10  instR3 (zll_rowround_rowround10_inR1[511:0], zll_rowround_rowround10_outR1);
  assign zll_columnround_columnround39_inR2 = zll_rowround_rowround10_outR1;
  ZLL_ColumnRound_columnround39  instR4 (zll_columnround_columnround39_inR2[511:0], zll_columnround_columnround39_outR2);
  assign zll_rowround_rowround10_inR2 = zll_columnround_columnround39_outR2;
  ZLL_RowRound_rowround10  instR5 (zll_rowround_rowround10_inR2[511:0], zll_rowround_rowround10_outR2);
  assign zll_columnround_columnround39_inR3 = zll_rowround_rowround10_outR2;
  ZLL_ColumnRound_columnround39  instR6 (zll_columnround_columnround39_inR3[511:0], zll_columnround_columnround39_outR3);
  assign zll_rowround_rowround10_inR3 = zll_columnround_columnround39_outR3;
  ZLL_RowRound_rowround10  instR7 (zll_rowround_rowround10_inR3[511:0], zll_rowround_rowround10_outR3);
  assign zll_columnround_columnround39_inR4 = zll_rowround_rowround10_outR3;
  ZLL_ColumnRound_columnround39  instR8 (zll_columnround_columnround39_inR4[511:0], zll_columnround_columnround39_outR4);
  assign zll_rowround_rowround10_inR4 = zll_columnround_columnround39_outR4;
  ZLL_RowRound_rowround10  instR9 (zll_rowround_rowround10_inR4[511:0], zll_rowround_rowround10_outR4);
  assign lit_in = zll_main_io_dr51_in[512:0];
  assign res = (lit_in[512] == 1'h0) ? {10'h201{1'h0}} : {1'h1, zll_rowround_rowround10_outR4};
endmodule

module ZLL_RowRound_rowround10 (input logic [511:0] arg0,
  output logic [511:0] res);
  logic [511:0] zll_rowround_rowround33_in;
  logic [511:0] zll_rowround_rowround9_in;
  logic [511:0] zll_rowround_rowround37_in;
  logic [511:0] zll_rowround_rowround25_in;
  logic [511:0] zll_rowround_rowround18_in;
  logic [511:0] zll_rowround_rowround35_in;
  logic [511:0] zll_rowround_rowround22_in;
  logic [511:0] zll_rowround_rowround4_in;
  logic [511:0] zll_rowround_rowround20_in;
  logic [511:0] zll_rowround_rowround19_in;
  logic [511:0] zll_rowround_rowround38_in;
  logic [511:0] zll_rowround_rowround5_in;
  logic [511:0] zll_rowround_rowround24_in;
  logic [127:0] zll_quarterround_quarterround15_in;
  logic [127:0] zll_quarterround_quarterround15_out;
  logic [511:0] zll_rowround_rowround15_in;
  logic [511:0] zll_rowround_rowround31_in;
  logic [511:0] zll_rowround_rowround1_in;
  logic [511:0] zll_rowround_rowround28_in;
  logic [127:0] zll_quarterround_quarterround15_inR1;
  logic [127:0] zll_quarterround_quarterround15_outR1;
  logic [511:0] zll_rowround_rowround39_in;
  logic [511:0] zll_rowround_rowround3_in;
  logic [511:0] zll_rowround_rowround12_in;
  logic [511:0] zll_rowround_rowround17_in;
  logic [511:0] zll_rowround_rowround32_in;
  logic [127:0] zll_quarterround_quarterround15_inR2;
  logic [127:0] zll_quarterround_quarterround15_outR2;
  logic [511:0] zll_rowround_rowround26_in;
  logic [511:0] zll_rowround_rowround11_in;
  logic [511:0] zll_rowround_rowround30_in;
  logic [511:0] zll_rowround_rowround8_in;
  logic [511:0] zll_rowround_rowround23_in;
  logic [127:0] zll_quarterround_quarterround15_inR3;
  logic [127:0] zll_quarterround_quarterround15_outR3;
  logic [511:0] zll_rowround_rowround34_in;
  logic [511:0] zll_rowround_rowround13_in;
  logic [511:0] zll_rowround_rowround_in;
  logic [511:0] zll_rowround_rowround2_in;
  logic [511:0] zll_rowround_rowround36_in;
  assign zll_rowround_rowround33_in = arg0;
  assign zll_rowround_rowround9_in = {zll_rowround_rowround33_in[479:448], zll_rowround_rowround33_in[511:480], zll_rowround_rowround33_in[447:416], zll_rowround_rowround33_in[415:384], zll_rowround_rowround33_in[383:352], zll_rowround_rowround33_in[351:320], zll_rowround_rowround33_in[319:288], zll_rowround_rowround33_in[287:256], zll_rowround_rowround33_in[255:224], zll_rowround_rowround33_in[223:192], zll_rowround_rowround33_in[191:160], zll_rowround_rowround33_in[159:128], zll_rowround_rowround33_in[127:96], zll_rowround_rowround33_in[95:64], zll_rowround_rowround33_in[63:32], zll_rowround_rowround33_in[31:0]};
  assign zll_rowround_rowround37_in = {zll_rowround_rowround9_in[447:416], zll_rowround_rowround9_in[511:480], zll_rowround_rowround9_in[479:448], zll_rowround_rowround9_in[415:384], zll_rowround_rowround9_in[383:352], zll_rowround_rowround9_in[351:320], zll_rowround_rowround9_in[319:288], zll_rowround_rowround9_in[287:256], zll_rowround_rowround9_in[255:224], zll_rowround_rowround9_in[223:192], zll_rowround_rowround9_in[191:160], zll_rowround_rowround9_in[159:128], zll_rowround_rowround9_in[127:96], zll_rowround_rowround9_in[95:64], zll_rowround_rowround9_in[63:32], zll_rowround_rowround9_in[31:0]};
  assign zll_rowround_rowround25_in = {zll_rowround_rowround37_in[511:480], zll_rowround_rowround37_in[383:352], zll_rowround_rowround37_in[479:448], zll_rowround_rowround37_in[447:416], zll_rowround_rowround37_in[415:384], zll_rowround_rowround37_in[351:320], zll_rowround_rowround37_in[319:288], zll_rowround_rowround37_in[287:256], zll_rowround_rowround37_in[255:224], zll_rowround_rowround37_in[223:192], zll_rowround_rowround37_in[191:160], zll_rowround_rowround37_in[159:128], zll_rowround_rowround37_in[127:96], zll_rowround_rowround37_in[95:64], zll_rowround_rowround37_in[63:32], zll_rowround_rowround37_in[31:0]};
  assign zll_rowround_rowround18_in = {zll_rowround_rowround25_in[511:480], zll_rowround_rowround25_in[479:448], zll_rowround_rowround25_in[351:320], zll_rowround_rowround25_in[447:416], zll_rowround_rowround25_in[415:384], zll_rowround_rowround25_in[383:352], zll_rowround_rowround25_in[319:288], zll_rowround_rowround25_in[287:256], zll_rowround_rowround25_in[255:224], zll_rowround_rowround25_in[223:192], zll_rowround_rowround25_in[191:160], zll_rowround_rowround25_in[159:128], zll_rowround_rowround25_in[127:96], zll_rowround_rowround25_in[95:64], zll_rowround_rowround25_in[63:32], zll_rowround_rowround25_in[31:0]};
  assign zll_rowround_rowround35_in = {zll_rowround_rowround18_in[511:480], zll_rowround_rowround18_in[479:448], zll_rowround_rowround18_in[287:256], zll_rowround_rowround18_in[447:416], zll_rowround_rowround18_in[415:384], zll_rowround_rowround18_in[383:352], zll_rowround_rowround18_in[351:320], zll_rowround_rowround18_in[319:288], zll_rowround_rowround18_in[255:224], zll_rowround_rowround18_in[223:192], zll_rowround_rowround18_in[191:160], zll_rowround_rowround18_in[159:128], zll_rowround_rowround18_in[127:96], zll_rowround_rowround18_in[95:64], zll_rowround_rowround18_in[63:32], zll_rowround_rowround18_in[31:0]};
  assign zll_rowround_rowround22_in = {zll_rowround_rowround35_in[511:480], zll_rowround_rowround35_in[479:448], zll_rowround_rowround35_in[447:416], zll_rowround_rowround35_in[415:384], zll_rowround_rowround35_in[383:352], zll_rowround_rowround35_in[351:320], zll_rowround_rowround35_in[255:224], zll_rowround_rowround35_in[319:288], zll_rowround_rowround35_in[287:256], zll_rowround_rowround35_in[223:192], zll_rowround_rowround35_in[191:160], zll_rowround_rowround35_in[159:128], zll_rowround_rowround35_in[127:96], zll_rowround_rowround35_in[95:64], zll_rowround_rowround35_in[63:32], zll_rowround_rowround35_in[31:0]};
  assign zll_rowround_rowround4_in = {zll_rowround_rowround22_in[511:480], zll_rowround_rowround22_in[479:448], zll_rowround_rowround22_in[447:416], zll_rowround_rowround22_in[415:384], zll_rowround_rowround22_in[383:352], zll_rowround_rowround22_in[351:320], zll_rowround_rowround22_in[223:192], zll_rowround_rowround22_in[319:288], zll_rowround_rowround22_in[287:256], zll_rowround_rowround22_in[255:224], zll_rowround_rowround22_in[191:160], zll_rowround_rowround22_in[159:128], zll_rowround_rowround22_in[127:96], zll_rowround_rowround22_in[95:64], zll_rowround_rowround22_in[63:32], zll_rowround_rowround22_in[31:0]};
  assign zll_rowround_rowround20_in = {zll_rowround_rowround4_in[511:480], zll_rowround_rowround4_in[479:448], zll_rowround_rowround4_in[447:416], zll_rowround_rowround4_in[415:384], zll_rowround_rowround4_in[383:352], zll_rowround_rowround4_in[351:320], zll_rowround_rowround4_in[319:288], zll_rowround_rowround4_in[287:256], zll_rowround_rowround4_in[255:224], zll_rowround_rowround4_in[191:160], zll_rowround_rowround4_in[223:192], zll_rowround_rowround4_in[159:128], zll_rowround_rowround4_in[127:96], zll_rowround_rowround4_in[95:64], zll_rowround_rowround4_in[63:32], zll_rowround_rowround4_in[31:0]};
  assign zll_rowround_rowround19_in = {zll_rowround_rowround20_in[511:480], zll_rowround_rowround20_in[479:448], zll_rowround_rowround20_in[447:416], zll_rowround_rowround20_in[415:384], zll_rowround_rowround20_in[383:352], zll_rowround_rowround20_in[351:320], zll_rowround_rowround20_in[319:288], zll_rowround_rowround20_in[287:256], zll_rowround_rowround20_in[255:224], zll_rowround_rowround20_in[159:128], zll_rowround_rowround20_in[223:192], zll_rowround_rowround20_in[191:160], zll_rowround_rowround20_in[127:96], zll_rowround_rowround20_in[95:64], zll_rowround_rowround20_in[63:32], zll_rowround_rowround20_in[31:0]};
  assign zll_rowround_rowround38_in = {zll_rowround_rowround19_in[511:480], zll_rowround_rowround19_in[127:96], zll_rowround_rowround19_in[479:448], zll_rowround_rowround19_in[447:416], zll_rowround_rowround19_in[415:384], zll_rowround_rowround19_in[383:352], zll_rowround_rowround19_in[351:320], zll_rowround_rowround19_in[319:288], zll_rowround_rowround19_in[287:256], zll_rowround_rowround19_in[255:224], zll_rowround_rowround19_in[223:192], zll_rowround_rowround19_in[191:160], zll_rowround_rowround19_in[159:128], zll_rowround_rowround19_in[95:64], zll_rowround_rowround19_in[63:32], zll_rowround_rowround19_in[31:0]};
  assign zll_rowround_rowround5_in = {zll_rowround_rowround38_in[511:480], zll_rowround_rowround38_in[479:448], zll_rowround_rowround38_in[95:64], zll_rowround_rowround38_in[447:416], zll_rowround_rowround38_in[415:384], zll_rowround_rowround38_in[383:352], zll_rowround_rowround38_in[351:320], zll_rowround_rowround38_in[319:288], zll_rowround_rowround38_in[287:256], zll_rowround_rowround38_in[255:224], zll_rowround_rowround38_in[223:192], zll_rowround_rowround38_in[191:160], zll_rowround_rowround38_in[159:128], zll_rowround_rowround38_in[127:96], zll_rowround_rowround38_in[63:32], zll_rowround_rowround38_in[31:0]};
  assign zll_rowround_rowround24_in = {zll_rowround_rowround5_in[511:480], zll_rowround_rowround5_in[479:448], zll_rowround_rowround5_in[447:416], zll_rowround_rowround5_in[415:384], zll_rowround_rowround5_in[383:352], zll_rowround_rowround5_in[351:320], zll_rowround_rowround5_in[63:32], zll_rowround_rowround5_in[319:288], zll_rowround_rowround5_in[287:256], zll_rowround_rowround5_in[255:224], zll_rowround_rowround5_in[223:192], zll_rowround_rowround5_in[191:160], zll_rowround_rowround5_in[159:128], zll_rowround_rowround5_in[127:96], zll_rowround_rowround5_in[95:64], zll_rowround_rowround5_in[31:0]};
  assign zll_quarterround_quarterround15_in = {zll_rowround_rowround24_in[255:224], zll_rowround_rowround24_in[287:256], zll_rowround_rowround24_in[511:480], zll_rowround_rowround24_in[159:128]};
  ZLL_QuarterRound_quarterround15  inst (zll_quarterround_quarterround15_in[127:0], zll_quarterround_quarterround15_out);
  assign zll_rowround_rowround15_in = {zll_rowround_rowround24_in[479:448], zll_rowround_rowround24_in[447:416], zll_rowround_rowround24_in[415:384], zll_rowround_rowround24_in[383:352], zll_rowround_rowround24_in[351:320], zll_rowround_rowround24_in[319:288], zll_rowround_rowround24_in[223:192], zll_rowround_rowround24_in[191:160], zll_rowround_rowround24_in[127:96], zll_rowround_rowround24_in[95:64], zll_rowround_rowround24_in[31:0], zll_rowround_rowround24_in[63:32], zll_quarterround_quarterround15_out};
  assign zll_rowround_rowround31_in = {zll_rowround_rowround15_in[511:480], zll_rowround_rowround15_in[479:448], zll_rowround_rowround15_in[447:416], zll_rowround_rowround15_in[415:384], zll_rowround_rowround15_in[383:352], zll_rowround_rowround15_in[351:320], zll_rowround_rowround15_in[319:288], zll_rowround_rowround15_in[287:256], zll_rowround_rowround15_in[255:224], zll_rowround_rowround15_in[223:192], zll_rowround_rowround15_in[191:160], zll_rowround_rowround15_in[159:128], zll_rowround_rowround15_in[127:0]};
  assign zll_rowround_rowround1_in = {zll_rowround_rowround31_in[511:480], zll_rowround_rowround31_in[479:448], zll_rowround_rowround31_in[447:416], zll_rowround_rowround31_in[415:384], zll_rowround_rowround31_in[383:352], zll_rowround_rowround31_in[351:320], zll_rowround_rowround31_in[127:96], zll_rowround_rowround31_in[319:288], zll_rowround_rowround31_in[287:256], zll_rowround_rowround31_in[255:224], zll_rowround_rowround31_in[223:192], zll_rowround_rowround31_in[191:160], zll_rowround_rowround31_in[159:128], zll_rowround_rowround31_in[95:64], zll_rowround_rowround31_in[63:32], zll_rowround_rowround31_in[31:0]};
  assign zll_rowround_rowround28_in = {zll_rowround_rowround1_in[511:480], zll_rowround_rowround1_in[479:448], zll_rowround_rowround1_in[63:32], zll_rowround_rowround1_in[447:416], zll_rowround_rowround1_in[415:384], zll_rowround_rowround1_in[383:352], zll_rowround_rowround1_in[351:320], zll_rowround_rowround1_in[319:288], zll_rowround_rowround1_in[287:256], zll_rowround_rowround1_in[255:224], zll_rowround_rowround1_in[223:192], zll_rowround_rowround1_in[191:160], zll_rowround_rowround1_in[159:128], zll_rowround_rowround1_in[127:96], zll_rowround_rowround1_in[95:64], zll_rowround_rowround1_in[31:0]};
  assign zll_quarterround_quarterround15_inR1 = {zll_rowround_rowround28_in[351:320], zll_rowround_rowround28_in[95:64], zll_rowround_rowround28_in[383:352], zll_rowround_rowround28_in[415:384]};
  ZLL_QuarterRound_quarterround15  instR1 (zll_quarterround_quarterround15_inR1[127:0], zll_quarterround_quarterround15_outR1);
  assign zll_rowround_rowround39_in = {zll_rowround_rowround28_in[511:480], zll_rowround_rowround28_in[479:448], zll_rowround_rowround28_in[447:416], zll_rowround_rowround28_in[319:288], zll_rowround_rowround28_in[287:256], zll_rowround_rowround28_in[255:224], zll_rowround_rowround28_in[31:0], zll_rowround_rowround28_in[223:192], zll_rowround_rowround28_in[191:160], zll_rowround_rowround28_in[159:128], zll_rowround_rowround28_in[127:96], zll_rowround_rowround28_in[63:32], zll_quarterround_quarterround15_outR1};
  assign zll_rowround_rowround3_in = {zll_rowround_rowround39_in[511:480], zll_rowround_rowround39_in[479:448], zll_rowround_rowround39_in[447:416], zll_rowround_rowround39_in[415:384], zll_rowround_rowround39_in[383:352], zll_rowround_rowround39_in[351:320], zll_rowround_rowround39_in[319:288], zll_rowround_rowround39_in[287:256], zll_rowround_rowround39_in[255:224], zll_rowround_rowround39_in[223:192], zll_rowround_rowround39_in[191:160], zll_rowround_rowround39_in[159:128], zll_rowround_rowround39_in[127:0]};
  assign zll_rowround_rowround12_in = {zll_rowround_rowround3_in[511:480], zll_rowround_rowround3_in[479:448], zll_rowround_rowround3_in[447:416], zll_rowround_rowround3_in[415:384], zll_rowround_rowround3_in[383:352], zll_rowround_rowround3_in[351:320], zll_rowround_rowround3_in[319:288], zll_rowround_rowround3_in[287:256], zll_rowround_rowround3_in[255:224], zll_rowround_rowround3_in[223:192], zll_rowround_rowround3_in[191:160], zll_rowround_rowround3_in[127:96], zll_rowround_rowround3_in[159:128], zll_rowround_rowround3_in[95:64], zll_rowround_rowround3_in[63:32], zll_rowround_rowround3_in[31:0]};
  assign zll_rowround_rowround17_in = {zll_rowround_rowround12_in[511:480], zll_rowround_rowround12_in[95:64], zll_rowround_rowround12_in[479:448], zll_rowround_rowround12_in[447:416], zll_rowround_rowround12_in[415:384], zll_rowround_rowround12_in[383:352], zll_rowround_rowround12_in[351:320], zll_rowround_rowround12_in[319:288], zll_rowround_rowround12_in[287:256], zll_rowround_rowround12_in[255:224], zll_rowround_rowround12_in[223:192], zll_rowround_rowround12_in[191:160], zll_rowround_rowround12_in[159:128], zll_rowround_rowround12_in[127:96], zll_rowround_rowround12_in[63:32], zll_rowround_rowround12_in[31:0]};
  assign zll_rowround_rowround32_in = {zll_rowround_rowround17_in[511:480], zll_rowround_rowround17_in[63:32], zll_rowround_rowround17_in[479:448], zll_rowround_rowround17_in[447:416], zll_rowround_rowround17_in[415:384], zll_rowround_rowround17_in[383:352], zll_rowround_rowround17_in[351:320], zll_rowround_rowround17_in[319:288], zll_rowround_rowround17_in[287:256], zll_rowround_rowround17_in[255:224], zll_rowround_rowround17_in[223:192], zll_rowround_rowround17_in[191:160], zll_rowround_rowround17_in[159:128], zll_rowround_rowround17_in[127:96], zll_rowround_rowround17_in[95:64], zll_rowround_rowround17_in[31:0]};
  assign zll_quarterround_quarterround15_inR2 = {zll_rowround_rowround32_in[159:128], zll_rowround_rowround32_in[191:160], zll_rowround_rowround32_in[223:192], zll_rowround_rowround32_in[287:256]};
  ZLL_QuarterRound_quarterround15  instR2 (zll_quarterround_quarterround15_inR2[127:0], zll_quarterround_quarterround15_outR2);
  assign zll_rowround_rowround26_in = {zll_rowround_rowround32_in[511:480], zll_rowround_rowround32_in[479:448], zll_rowround_rowround32_in[447:416], zll_rowround_rowround32_in[415:384], zll_rowround_rowround32_in[383:352], zll_rowround_rowround32_in[351:320], zll_rowround_rowround32_in[319:288], zll_rowround_rowround32_in[255:224], zll_rowround_rowround32_in[127:96], zll_rowround_rowround32_in[31:0], zll_rowround_rowround32_in[95:64], zll_rowround_rowround32_in[63:32], zll_quarterround_quarterround15_outR2};
  assign zll_rowround_rowround11_in = {zll_rowround_rowround26_in[511:480], zll_rowround_rowround26_in[479:448], zll_rowround_rowround26_in[447:416], zll_rowround_rowround26_in[415:384], zll_rowround_rowround26_in[383:352], zll_rowround_rowround26_in[351:320], zll_rowround_rowround26_in[319:288], zll_rowround_rowround26_in[287:256], zll_rowround_rowround26_in[255:224], zll_rowround_rowround26_in[223:192], zll_rowround_rowround26_in[191:160], zll_rowround_rowround26_in[159:128], zll_rowround_rowround26_in[127:0]};
  assign zll_rowround_rowround30_in = {zll_rowround_rowround11_in[511:480], zll_rowround_rowround11_in[479:448], zll_rowround_rowround11_in[447:416], zll_rowround_rowround11_in[415:384], zll_rowround_rowround11_in[383:352], zll_rowround_rowround11_in[351:320], zll_rowround_rowround11_in[319:288], zll_rowround_rowround11_in[287:256], zll_rowround_rowround11_in[127:96], zll_rowround_rowround11_in[255:224], zll_rowround_rowround11_in[223:192], zll_rowround_rowround11_in[191:160], zll_rowround_rowround11_in[159:128], zll_rowround_rowround11_in[95:64], zll_rowround_rowround11_in[63:32], zll_rowround_rowround11_in[31:0]};
  assign zll_rowround_rowround8_in = {zll_rowround_rowround30_in[511:480], zll_rowround_rowround30_in[479:448], zll_rowround_rowround30_in[447:416], zll_rowround_rowround30_in[415:384], zll_rowround_rowround30_in[383:352], zll_rowround_rowround30_in[351:320], zll_rowround_rowround30_in[319:288], zll_rowround_rowround30_in[287:256], zll_rowround_rowround30_in[255:224], zll_rowround_rowround30_in[95:64], zll_rowround_rowround30_in[223:192], zll_rowround_rowround30_in[191:160], zll_rowround_rowround30_in[159:128], zll_rowround_rowround30_in[127:96], zll_rowround_rowround30_in[63:32], zll_rowround_rowround30_in[31:0]};
  assign zll_rowround_rowround23_in = {zll_rowround_rowround8_in[511:480], zll_rowround_rowround8_in[479:448], zll_rowround_rowround8_in[447:416], zll_rowround_rowround8_in[415:384], zll_rowround_rowround8_in[383:352], zll_rowround_rowround8_in[63:32], zll_rowround_rowround8_in[351:320], zll_rowround_rowround8_in[319:288], zll_rowround_rowround8_in[287:256], zll_rowround_rowround8_in[255:224], zll_rowround_rowround8_in[223:192], zll_rowround_rowround8_in[191:160], zll_rowround_rowround8_in[159:128], zll_rowround_rowround8_in[127:96], zll_rowround_rowround8_in[95:64], zll_rowround_rowround8_in[31:0]};
  assign zll_quarterround_quarterround15_inR3 = {zll_rowround_rowround23_in[159:128], zll_rowround_rowround23_in[511:480], zll_rowround_rowround23_in[415:384], zll_rowround_rowround23_in[319:288]};
  ZLL_QuarterRound_quarterround15  instR3 (zll_quarterround_quarterround15_inR3[127:0], zll_quarterround_quarterround15_outR3);
  assign zll_rowround_rowround34_in = {zll_rowround_rowround23_in[479:448], zll_rowround_rowround23_in[447:416], zll_rowround_rowround23_in[383:352], zll_rowround_rowround23_in[31:0], zll_rowround_rowround23_in[351:320], zll_rowround_rowround23_in[287:256], zll_rowround_rowround23_in[255:224], zll_rowround_rowround23_in[223:192], zll_rowround_rowround23_in[191:160], zll_rowround_rowround23_in[127:96], zll_rowround_rowround23_in[95:64], zll_rowround_rowround23_in[63:32], zll_quarterround_quarterround15_outR3};
  assign zll_rowround_rowround13_in = {zll_rowround_rowround34_in[511:480], zll_rowround_rowround34_in[479:448], zll_rowround_rowround34_in[447:416], zll_rowround_rowround34_in[415:384], zll_rowround_rowround34_in[383:352], zll_rowround_rowround34_in[351:320], zll_rowround_rowround34_in[319:288], zll_rowround_rowround34_in[287:256], zll_rowround_rowround34_in[255:224], zll_rowround_rowround34_in[223:192], zll_rowround_rowround34_in[191:160], zll_rowround_rowround34_in[159:128], zll_rowround_rowround34_in[127:0]};
  assign zll_rowround_rowround_in = {zll_rowround_rowround13_in[511:480], zll_rowround_rowround13_in[479:448], zll_rowround_rowround13_in[447:416], zll_rowround_rowround13_in[415:384], zll_rowround_rowround13_in[383:352], zll_rowround_rowround13_in[351:320], zll_rowround_rowround13_in[319:288], zll_rowround_rowround13_in[127:96], zll_rowround_rowround13_in[287:256], zll_rowround_rowround13_in[255:224], zll_rowround_rowround13_in[223:192], zll_rowround_rowround13_in[191:160], zll_rowround_rowround13_in[159:128], zll_rowround_rowround13_in[95:64], zll_rowround_rowround13_in[63:32], zll_rowround_rowround13_in[31:0]};
  assign zll_rowround_rowround2_in = {zll_rowround_rowround_in[95:64], zll_rowround_rowround_in[511:480], zll_rowround_rowround_in[479:448], zll_rowround_rowround_in[447:416], zll_rowround_rowround_in[415:384], zll_rowround_rowround_in[383:352], zll_rowround_rowround_in[351:320], zll_rowround_rowround_in[319:288], zll_rowround_rowround_in[287:256], zll_rowround_rowround_in[255:224], zll_rowround_rowround_in[223:192], zll_rowround_rowround_in[191:160], zll_rowround_rowround_in[159:128], zll_rowround_rowround_in[127:96], zll_rowround_rowround_in[63:32], zll_rowround_rowround_in[31:0]};
  assign zll_rowround_rowround36_in = {zll_rowround_rowround2_in[511:480], zll_rowround_rowround2_in[479:448], zll_rowround_rowround2_in[447:416], zll_rowround_rowround2_in[415:384], zll_rowround_rowround2_in[383:352], zll_rowround_rowround2_in[351:320], zll_rowround_rowround2_in[319:288], zll_rowround_rowround2_in[287:256], zll_rowround_rowround2_in[255:224], zll_rowround_rowround2_in[63:32], zll_rowround_rowround2_in[223:192], zll_rowround_rowround2_in[191:160], zll_rowround_rowround2_in[159:128], zll_rowround_rowround2_in[127:96], zll_rowround_rowround2_in[95:64], zll_rowround_rowround2_in[31:0]};
  assign res = {zll_rowround_rowround36_in[319:288], zll_rowround_rowround36_in[63:32], zll_rowround_rowround36_in[415:384], zll_rowround_rowround36_in[287:256], zll_rowround_rowround36_in[127:96], zll_rowround_rowround36_in[95:64], zll_rowround_rowround36_in[447:416], zll_rowround_rowround36_in[479:448], zll_rowround_rowround36_in[351:320], zll_rowround_rowround36_in[383:352], zll_rowround_rowround36_in[191:160], zll_rowround_rowround36_in[159:128], zll_rowround_rowround36_in[511:480], zll_rowround_rowround36_in[223:192], zll_rowround_rowround36_in[31:0], zll_rowround_rowround36_in[255:224]};
endmodule

module ZLL_Main_out2 (input logic [1025:0] arg0,
  output logic [512:0] res);
  logic [1025:0] zll_main_out21_in;
  assign zll_main_out21_in = arg0;
  assign res = zll_main_out21_in[512:0];
endmodule